// DE2_115_SOPC.v

// Generated using ACDS version 13.1 182 at 2015.03.26.09:07:03

`timescale 1 ps / 1 ps
module DE2_115_SOPC (
		input  wire        clk_50_clk,                                                    //                            clk_50.clk
		input  wire        reset_reset_n,                                                 //                             reset.reset_n
		output wire [10:0] sdram_wire_addr,                                               //                        sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                                 //                                  .ba
		output wire        sdram_wire_cas_n,                                              //                                  .cas_n
		output wire        sdram_wire_cke,                                                //                                  .cke
		output wire        sdram_wire_cs_n,                                               //                                  .cs_n
		inout  wire [31:0] sdram_wire_dq,                                                 //                                  .dq
		output wire [3:0]  sdram_wire_dqm,                                                //                                  .dqm
		output wire        sdram_wire_ras_n,                                              //                                  .ras_n
		output wire        sdram_wire_we_n,                                               //                                  .we_n
		inout  wire [15:0] sram_conduit_end_DQ,                                           //                  sram_conduit_end.DQ
		output wire [19:0] sram_conduit_end_ADDR,                                         //                                  .ADDR
		output wire        sram_conduit_end_UB_n,                                         //                                  .UB_n
		output wire        sram_conduit_end_LB_n,                                         //                                  .LB_n
		output wire        sram_conduit_end_WE_n,                                         //                                  .WE_n
		output wire        sram_conduit_end_CE_n,                                         //                                  .CE_n
		output wire        sram_conduit_end_OE_n,                                         //                                  .OE_n
		output wire [22:0] tristate_conduit_bridge_flash_out_address_to_the_cfi_flash,    // tristate_conduit_bridge_flash_out.address_to_the_cfi_flash
		inout  wire [7:0]  tristate_conduit_bridge_flash_out_tri_state_bridge_flash_data, //                                  .tri_state_bridge_flash_data
		output wire [0:0]  tristate_conduit_bridge_flash_out_write_n_to_the_cfi_flash,    //                                  .write_n_to_the_cfi_flash
		output wire [0:0]  tristate_conduit_bridge_flash_out_select_n_to_the_cfi_flash,   //                                  .select_n_to_the_cfi_flash
		output wire [0:0]  tristate_conduit_bridge_flash_out_read_n_to_the_cfi_flash,     //                                  .read_n_to_the_cfi_flash
		output wire        altpll_sdram_clk,                                              //                      altpll_sdram.clk
		output wire        altpll_25_clk,                                                 //                         altpll_25.clk
		input  wire        pll_areset_conduit_export,                                     //                pll_areset_conduit.export
		output wire        pll_locked_conduit_export,                                     //                pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export,                                  //             pll_phasedone_conduit.export
		output wire        altpll_sys_clk,                                                //                        altpll_sys.clk
		output wire        altpll_io_clk,                                                 //                         altpll_io.clk
		input  wire [3:0]  key_external_connection_export,                                //           key_external_connection.export
		input  wire [17:0] sw_external_connection_export,                                 //            sw_external_connection.export
		output wire [8:0]  ledg_external_connection_export,                               //          ledg_external_connection.export
		output wire [17:0] ledr_external_connection_export,                               //          ledr_external_connection.export
		input  wire        rs232_external_connection_rxd,                                 //         rs232_external_connection.rxd
		output wire        rs232_external_connection_txd,                                 //                                  .txd
		input  wire        rs232_external_connection_cts_n,                               //                                  .cts_n
		output wire        rs232_external_connection_rts_n,                               //                                  .rts_n
		output wire        i2c_scl_external_connection_export,                            //       i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export,                            //       i2c_sda_external_connection.export
		output wire        eep_i2c_scl_external_connection_export,                        //   eep_i2c_scl_external_connection.export
		inout  wire        eep_i2c_sda_external_connection_export,                        //   eep_i2c_sda_external_connection.export
		output wire        lcd_external_RS,                                               //                      lcd_external.RS
		output wire        lcd_external_RW,                                               //                                  .RW
		inout  wire [7:0]  lcd_external_data,                                             //                                  .data
		output wire        lcd_external_E,                                                //                                  .E
		input  wire        ir_external_connection_export,                                 //            ir_external_connection.export
		output wire        sd_clk_external_connection_export,                             //        sd_clk_external_connection.export
		inout  wire        sd_cmd_external_connection_export,                             //        sd_cmd_external_connection.export
		inout  wire [3:0]  sd_dat_external_connection_export,                             //        sd_dat_external_connection.export
		input  wire        sd_wp_n_external_connection_export,                            //       sd_wp_n_external_connection.export
		output wire [63:0] seg7_conduit_end_export,                                       //                  seg7_conduit_end.export
		input  wire        sma_in_external_connection_export,                             //        sma_in_external_connection.export
		output wire        sma_out_external_connection_export,                            //       sma_out_external_connection.export
		output wire        audio_conduit_end_XCK,                                         //                 audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                                      //                                  .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                                      //                                  .ADCLRC
		output wire        audio_conduit_end_DACDAT,                                      //                                  .DACDAT
		input  wire        audio_conduit_end_DACLRC,                                      //                                  .DACLRC
		input  wire        audio_conduit_end_BCLK,                                        //                                  .BCLK
		inout  wire [15:0] usb_conduit_end_DATA,                                          //                   usb_conduit_end.DATA
		output wire [1:0]  usb_conduit_end_ADDR,                                          //                                  .ADDR
		output wire        usb_conduit_end_RD_N,                                          //                                  .RD_N
		output wire        usb_conduit_end_WR_N,                                          //                                  .WR_N
		output wire        usb_conduit_end_CS_N,                                          //                                  .CS_N
		output wire        usb_conduit_end_RST_N,                                         //                                  .RST_N
		input  wire        usb_conduit_end_INT0,                                          //                                  .INT0
		input  wire        usb_conduit_end_INT1,                                          //                                  .INT1
		output wire        can_top_0_conduit_end_tx_o,                                    //             can_top_0_conduit_end.tx_o
		input  wire        can_top_0_conduit_end_rx_i,                                    //                                  .rx_i
		output wire        can_top_0_conduit_end_clkout_o,                                //                                  .clkout_o
		output wire        can_top_0_conduit_end_bus_off_on,                              //                                  .bus_off_on
		input  wire        uart_0_external_connection_rxd,                                //        uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd,                                //                                  .txd
		input  wire        uart_1_external_connection_rxd,                                //        uart_1_external_connection.rxd
		output wire        uart_1_external_connection_txd,                                //                                  .txd
		input  wire        tse_pcs_mac_tx_clock_connection_clk,                           //   tse_pcs_mac_tx_clock_connection.clk
		input  wire        tse_pcs_mac_rx_clock_connection_clk,                           //   tse_pcs_mac_rx_clock_connection.clk
		input  wire        tse_mac_status_connection_set_10,                              //         tse_mac_status_connection.set_10
		input  wire        tse_mac_status_connection_set_1000,                            //                                  .set_1000
		output wire        tse_mac_status_connection_eth_mode,                            //                                  .eth_mode
		output wire        tse_mac_status_connection_ena_10,                              //                                  .ena_10
		input  wire [3:0]  tse_mac_rgmii_connection_rgmii_in,                             //          tse_mac_rgmii_connection.rgmii_in
		output wire [3:0]  tse_mac_rgmii_connection_rgmii_out,                            //                                  .rgmii_out
		input  wire        tse_mac_rgmii_connection_rx_control,                           //                                  .rx_control
		output wire        tse_mac_rgmii_connection_tx_control,                           //                                  .tx_control
		output wire        tse_mac_mdio_connection_mdc,                                   //           tse_mac_mdio_connection.mdc
		input  wire        tse_mac_mdio_connection_mdio_in,                               //                                  .mdio_in
		output wire        tse_mac_mdio_connection_mdio_out,                              //                                  .mdio_out
		output wire        tse_mac_mdio_connection_mdio_oen,                              //                                  .mdio_oen
		input  wire        tse_mac_misc_connection_ff_tx_crc_fwd,                         //           tse_mac_misc_connection.ff_tx_crc_fwd
		output wire        tse_mac_misc_connection_ff_tx_septy,                           //                                  .ff_tx_septy
		output wire        tse_mac_misc_connection_tx_ff_uflow,                           //                                  .tx_ff_uflow
		output wire        tse_mac_misc_connection_ff_tx_a_full,                          //                                  .ff_tx_a_full
		output wire        tse_mac_misc_connection_ff_tx_a_empty,                         //                                  .ff_tx_a_empty
		output wire [17:0] tse_mac_misc_connection_rx_err_stat,                           //                                  .rx_err_stat
		output wire [3:0]  tse_mac_misc_connection_rx_frm_type,                           //                                  .rx_frm_type
		output wire        tse_mac_misc_connection_ff_rx_dsav,                            //                                  .ff_rx_dsav
		output wire        tse_mac_misc_connection_ff_rx_a_full,                          //                                  .ff_rx_a_full
		output wire        tse_mac_misc_connection_ff_rx_a_empty                          //                                  .ff_rx_a_empty
	);

	wire         vic_0_interrupt_controller_out_valid;                                    // vic_0:interrupt_controller_out_valid -> cpu:eic_port_valid
	wire  [44:0] vic_0_interrupt_controller_out_data;                                     // vic_0:interrupt_controller_out_data -> cpu:eic_port_data
	wire   [7:0] tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_in;    // tristate_conduit_bridge_flash:tcs_tri_state_bridge_flash_data_in -> tristate_conduit_pin_sharer_flash:tri_state_bridge_flash_data_in
	wire   [7:0] tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_out;   // tristate_conduit_pin_sharer_flash:tri_state_bridge_flash_data -> tristate_conduit_bridge_flash:tcs_tri_state_bridge_flash_data
	wire         tristate_conduit_pin_sharer_flash_tcm_grant;                             // tristate_conduit_bridge_flash:grant -> tristate_conduit_pin_sharer_flash:grant
	wire   [0:0] tristate_conduit_pin_sharer_flash_tcm_select_n_to_the_cfi_flash_out;     // tristate_conduit_pin_sharer_flash:select_n_to_the_cfi_flash -> tristate_conduit_bridge_flash:tcs_select_n_to_the_cfi_flash
	wire         tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_outen; // tristate_conduit_pin_sharer_flash:tri_state_bridge_flash_data_outen -> tristate_conduit_bridge_flash:tcs_tri_state_bridge_flash_data_outen
	wire         tristate_conduit_pin_sharer_flash_tcm_request;                           // tristate_conduit_pin_sharer_flash:request -> tristate_conduit_bridge_flash:request
	wire   [0:0] tristate_conduit_pin_sharer_flash_tcm_write_n_to_the_cfi_flash_out;      // tristate_conduit_pin_sharer_flash:write_n_to_the_cfi_flash -> tristate_conduit_bridge_flash:tcs_write_n_to_the_cfi_flash
	wire   [0:0] tristate_conduit_pin_sharer_flash_tcm_read_n_to_the_cfi_flash_out;       // tristate_conduit_pin_sharer_flash:read_n_to_the_cfi_flash -> tristate_conduit_bridge_flash:tcs_read_n_to_the_cfi_flash
	wire  [22:0] tristate_conduit_pin_sharer_flash_tcm_address_to_the_cfi_flash_out;      // tristate_conduit_pin_sharer_flash:address_to_the_cfi_flash -> tristate_conduit_bridge_flash:tcs_address_to_the_cfi_flash
	wire         cfi_flash_tcm_chipselect_n_out;                                          // cfi_flash:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_flash:tcs0_chipselect_n_out
	wire         cfi_flash_tcm_grant;                                                     // tristate_conduit_pin_sharer_flash:tcs0_grant -> cfi_flash:tcm_grant
	wire         cfi_flash_tcm_data_outen;                                                // cfi_flash:tcm_data_outen -> tristate_conduit_pin_sharer_flash:tcs0_data_outen
	wire         cfi_flash_tcm_request;                                                   // cfi_flash:tcm_request -> tristate_conduit_pin_sharer_flash:tcs0_request
	wire   [7:0] cfi_flash_tcm_data_out;                                                  // cfi_flash:tcm_data_out -> tristate_conduit_pin_sharer_flash:tcs0_data_out
	wire         cfi_flash_tcm_write_n_out;                                               // cfi_flash:tcm_write_n_out -> tristate_conduit_pin_sharer_flash:tcs0_write_n_out
	wire  [22:0] cfi_flash_tcm_address_out;                                               // cfi_flash:tcm_address_out -> tristate_conduit_pin_sharer_flash:tcs0_address_out
	wire   [7:0] cfi_flash_tcm_data_in;                                                   // tristate_conduit_pin_sharer_flash:tcs0_data_in -> cfi_flash:tcm_data_in
	wire         cfi_flash_tcm_read_n_out;                                                // cfi_flash:tcm_read_n_out -> tristate_conduit_pin_sharer_flash:tcs0_read_n_out
	wire         sgdma_tx_out_endofpacket;                                                // sgdma_tx:out_endofpacket -> tse:ff_tx_eop
	wire         sgdma_tx_out_valid;                                                      // sgdma_tx:out_valid -> tse:ff_tx_wren
	wire         sgdma_tx_out_startofpacket;                                              // sgdma_tx:out_startofpacket -> tse:ff_tx_sop
	wire         sgdma_tx_out_error;                                                      // sgdma_tx:out_error -> tse:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                                      // sgdma_tx:out_empty -> tse:ff_tx_mod
	wire  [31:0] sgdma_tx_out_data;                                                       // sgdma_tx:out_data -> tse:ff_tx_data
	wire         sgdma_tx_out_ready;                                                      // tse:ff_tx_rdy -> sgdma_tx:out_ready
	wire         mm_interconnect_0_tse_control_port_waitrequest;                          // tse:waitrequest -> mm_interconnect_0:tse_control_port_waitrequest
	wire  [31:0] mm_interconnect_0_tse_control_port_writedata;                            // mm_interconnect_0:tse_control_port_writedata -> tse:writedata
	wire   [7:0] mm_interconnect_0_tse_control_port_address;                              // mm_interconnect_0:tse_control_port_address -> tse:address
	wire         mm_interconnect_0_tse_control_port_write;                                // mm_interconnect_0:tse_control_port_write -> tse:write
	wire         mm_interconnect_0_tse_control_port_read;                                 // mm_interconnect_0:tse_control_port_read -> tse:read
	wire  [31:0] mm_interconnect_0_tse_control_port_readdata;                             // tse:readdata -> mm_interconnect_0:tse_control_port_readdata
	wire  [31:0] mm_interconnect_0_vic_0_csr_access_writedata;                            // mm_interconnect_0:vic_0_csr_access_writedata -> vic_0:csr_access_writedata
	wire   [7:0] mm_interconnect_0_vic_0_csr_access_address;                              // mm_interconnect_0:vic_0_csr_access_address -> vic_0:csr_access_address
	wire         mm_interconnect_0_vic_0_csr_access_write;                                // mm_interconnect_0:vic_0_csr_access_write -> vic_0:csr_access_write
	wire         mm_interconnect_0_vic_0_csr_access_read;                                 // mm_interconnect_0:vic_0_csr_access_read -> vic_0:csr_access_read
	wire  [31:0] mm_interconnect_0_vic_0_csr_access_readdata;                             // vic_0:csr_access_readdata -> mm_interconnect_0:vic_0_csr_access_readdata
	wire         sgdma_rx_m_write_waitrequest;                                            // mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_writedata;                                              // sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	wire  [31:0] sgdma_rx_m_write_address;                                                // sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	wire         sgdma_rx_m_write_write;                                                  // sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	wire   [3:0] sgdma_rx_m_write_byteenable;                                             // sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                     // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                       // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                         // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                           // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                            // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                        // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                     // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                      // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cfi_flash_uas_waitrequest;                             // cfi_flash:uas_waitrequest -> mm_interconnect_0:cfi_flash_uas_waitrequest
	wire   [0:0] mm_interconnect_0_cfi_flash_uas_burstcount;                              // mm_interconnect_0:cfi_flash_uas_burstcount -> cfi_flash:uas_burstcount
	wire   [7:0] mm_interconnect_0_cfi_flash_uas_writedata;                               // mm_interconnect_0:cfi_flash_uas_writedata -> cfi_flash:uas_writedata
	wire  [22:0] mm_interconnect_0_cfi_flash_uas_address;                                 // mm_interconnect_0:cfi_flash_uas_address -> cfi_flash:uas_address
	wire         mm_interconnect_0_cfi_flash_uas_lock;                                    // mm_interconnect_0:cfi_flash_uas_lock -> cfi_flash:uas_lock
	wire         mm_interconnect_0_cfi_flash_uas_write;                                   // mm_interconnect_0:cfi_flash_uas_write -> cfi_flash:uas_write
	wire         mm_interconnect_0_cfi_flash_uas_read;                                    // mm_interconnect_0:cfi_flash_uas_read -> cfi_flash:uas_read
	wire   [7:0] mm_interconnect_0_cfi_flash_uas_readdata;                                // cfi_flash:uas_readdata -> mm_interconnect_0:cfi_flash_uas_readdata
	wire         mm_interconnect_0_cfi_flash_uas_debugaccess;                             // mm_interconnect_0:cfi_flash_uas_debugaccess -> cfi_flash:uas_debugaccess
	wire         mm_interconnect_0_cfi_flash_uas_readdatavalid;                           // cfi_flash:uas_readdatavalid -> mm_interconnect_0:cfi_flash_uas_readdatavalid
	wire   [0:0] mm_interconnect_0_cfi_flash_uas_byteenable;                              // mm_interconnect_0:cfi_flash_uas_byteenable -> cfi_flash:uas_byteenable
	wire         sgdma_tx_descriptor_read_waitrequest;                                    // mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                                        // sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                                           // sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                                       // mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_readdatavalid;                                  // mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                                // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                                  // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                               // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire         mm_interconnect_0_sgdma_tx_csr_write;                                    // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire         mm_interconnect_0_sgdma_tx_csr_read;                                     // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                                 // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire  [15:0] mm_interconnect_0_uart_1_s1_writedata;                                   // mm_interconnect_0:uart_1_s1_writedata -> uart_1:writedata
	wire   [2:0] mm_interconnect_0_uart_1_s1_address;                                     // mm_interconnect_0:uart_1_s1_address -> uart_1:address
	wire         mm_interconnect_0_uart_1_s1_chipselect;                                  // mm_interconnect_0:uart_1_s1_chipselect -> uart_1:chipselect
	wire         mm_interconnect_0_uart_1_s1_write;                                       // mm_interconnect_0:uart_1_s1_write -> uart_1:write_n
	wire         mm_interconnect_0_uart_1_s1_read;                                        // mm_interconnect_0:uart_1_s1_read -> uart_1:read_n
	wire  [15:0] mm_interconnect_0_uart_1_s1_readdata;                                    // uart_1:readdata -> mm_interconnect_0:uart_1_s1_readdata
	wire         mm_interconnect_0_uart_1_s1_begintransfer;                               // mm_interconnect_0:uart_1_s1_begintransfer -> uart_1:begintransfer
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                      // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                       // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                        // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire  [10:0] mm_interconnect_0_clock_crossing_io_s0_address;                          // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                            // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                             // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                         // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                      // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                    // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                       // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         sgdma_rx_descriptor_read_waitrequest;                                    // mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                                        // sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                                           // sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                                       // mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_readdatavalid;                                  // mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire  [31:0] mm_interconnect_0_sma_out_s1_writedata;                                  // mm_interconnect_0:sma_out_s1_writedata -> sma_out:writedata
	wire   [1:0] mm_interconnect_0_sma_out_s1_address;                                    // mm_interconnect_0:sma_out_s1_address -> sma_out:address
	wire         mm_interconnect_0_sma_out_s1_chipselect;                                 // mm_interconnect_0:sma_out_s1_chipselect -> sma_out:chipselect
	wire         mm_interconnect_0_sma_out_s1_write;                                      // mm_interconnect_0:sma_out_s1_write -> sma_out:write_n
	wire  [31:0] mm_interconnect_0_sma_out_s1_readdata;                                   // sma_out:readdata -> mm_interconnect_0:sma_out_s1_readdata
	wire         sgdma_rx_descriptor_write_waitrequest;                                   // mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                                     // sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	wire  [31:0] sgdma_rx_descriptor_write_address;                                       // sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                                         // sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	wire   [3:0] cpu_instruction_master_burstcount;                                       // cpu:i_burstcount -> mm_interconnect_0:cpu_instruction_master_burstcount
	wire         cpu_instruction_master_waitrequest;                                      // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                          // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                             // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                         // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                                    // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [15:0] mm_interconnect_0_usb_hc_writedata;                                      // mm_interconnect_0:usb_hc_writedata -> usb:avs_hc_writedata_iDATA
	wire   [0:0] mm_interconnect_0_usb_hc_address;                                        // mm_interconnect_0:usb_hc_address -> usb:avs_hc_address_iADDR
	wire         mm_interconnect_0_usb_hc_chipselect;                                     // mm_interconnect_0:usb_hc_chipselect -> usb:avs_hc_chipselect_n_iCS_N
	wire         mm_interconnect_0_usb_hc_write;                                          // mm_interconnect_0:usb_hc_write -> usb:avs_hc_write_n_iWR_N
	wire         mm_interconnect_0_usb_hc_read;                                           // mm_interconnect_0:usb_hc_read -> usb:avs_hc_read_n_iRD_N
	wire  [15:0] mm_interconnect_0_usb_hc_readdata;                                       // usb:avs_hc_readdata_oDATA -> mm_interconnect_0:usb_hc_readdata
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;                        // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire   [9:0] mm_interconnect_0_descriptor_memory_s1_address;                          // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;                       // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire         mm_interconnect_0_descriptor_memory_s1_clken;                            // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_0_descriptor_memory_s1_write;                            // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;                         // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;                       // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire   [1:0] mm_interconnect_0_sma_in_s1_address;                                     // mm_interconnect_0:sma_in_s1_address -> sma_in:address
	wire  [31:0] mm_interconnect_0_sma_in_s1_readdata;                                    // sma_in:readdata -> mm_interconnect_0:sma_in_s1_readdata
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                           // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                             // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                          // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                               // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_onchip_memory2_s1_write;                               // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                            // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                          // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                                // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                                  // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                               // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire         mm_interconnect_0_sgdma_rx_csr_write;                                    // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire         mm_interconnect_0_sgdma_rx_csr_read;                                     // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                                 // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_writedata;                           // mm_interconnect_0:sram_avalon_slave_writedata -> sram:s_writedata
	wire  [19:0] mm_interconnect_0_sram_avalon_slave_address;                             // mm_interconnect_0:sram_avalon_slave_address -> sram:s_address
	wire         mm_interconnect_0_sram_avalon_slave_chipselect;                          // mm_interconnect_0:sram_avalon_slave_chipselect -> sram:s_chipselect_n
	wire         mm_interconnect_0_sram_avalon_slave_write;                               // mm_interconnect_0:sram_avalon_slave_write -> sram:s_write_n
	wire         mm_interconnect_0_sram_avalon_slave_read;                                // mm_interconnect_0:sram_avalon_slave_read -> sram:s_read_n
	wire  [15:0] mm_interconnect_0_sram_avalon_slave_readdata;                            // sram:s_readdata -> mm_interconnect_0:sram_avalon_slave_readdata
	wire   [1:0] mm_interconnect_0_sram_avalon_slave_byteenable;                          // mm_interconnect_0:sram_avalon_slave_byteenable -> sram:s_byteenable_n
	wire  [15:0] mm_interconnect_0_usb_dc_writedata;                                      // mm_interconnect_0:usb_dc_writedata -> usb:avs_dc_writedata_iDATA
	wire   [0:0] mm_interconnect_0_usb_dc_address;                                        // mm_interconnect_0:usb_dc_address -> usb:avs_dc_address_iADDR
	wire         mm_interconnect_0_usb_dc_chipselect;                                     // mm_interconnect_0:usb_dc_chipselect -> usb:avs_dc_chipselect_n_iCS_N
	wire         mm_interconnect_0_usb_dc_write;                                          // mm_interconnect_0:usb_dc_write -> usb:avs_dc_write_n_iWR_N
	wire         mm_interconnect_0_usb_dc_read;                                           // mm_interconnect_0:usb_dc_read -> usb:avs_dc_read_n_iRD_N
	wire  [15:0] mm_interconnect_0_usb_dc_readdata;                                       // usb:avs_dc_readdata_oDATA -> mm_interconnect_0:usb_dc_readdata
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                   // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                     // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_chipselect;                                  // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire         mm_interconnect_0_uart_0_s1_write;                                       // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire         mm_interconnect_0_uart_0_s1_read;                                        // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                    // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                               // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                  // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                    // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [22:0] mm_interconnect_0_sdram_s1_address;                                      // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                   // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                        // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                         // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                     // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                   // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_writedata;                          // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire   [2:0] mm_interconnect_0_audio_avalon_slave_address;                            // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire         mm_interconnect_0_audio_avalon_slave_write;                              // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire         mm_interconnect_0_audio_avalon_slave_read;                               // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire  [15:0] mm_interconnect_0_audio_avalon_slave_readdata;                           // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire         cpu_data_master_waitrequest;                                             // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                               // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                                 // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                                   // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                                    // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                                // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                             // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                              // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         sgdma_tx_descriptor_write_waitrequest;                                   // mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                                     // sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	wire  [31:0] sgdma_tx_descriptor_write_address;                                       // sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                                         // sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	wire  [31:0] mm_interconnect_0_can_top_0_avalon_slave_0_writedata;                    // mm_interconnect_0:can_top_0_avalon_slave_0_writedata -> can_top_0:av_dat_i
	wire   [7:0] mm_interconnect_0_can_top_0_avalon_slave_0_address;                      // mm_interconnect_0:can_top_0_avalon_slave_0_address -> can_top_0:av_adr_i
	wire         mm_interconnect_0_can_top_0_avalon_slave_0_chipselect;                   // mm_interconnect_0:can_top_0_avalon_slave_0_chipselect -> can_top_0:av_cs_i
	wire         mm_interconnect_0_can_top_0_avalon_slave_0_write;                        // mm_interconnect_0:can_top_0_avalon_slave_0_write -> can_top_0:av_wr_i
	wire  [31:0] mm_interconnect_0_can_top_0_avalon_slave_0_readdata;                     // can_top_0:av_dat_o -> mm_interconnect_0:can_top_0_avalon_slave_0_readdata
	wire         sgdma_tx_m_read_waitrequest;                                             // mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                                 // sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                                    // sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	wire  [31:0] sgdma_tx_m_read_readdata;                                                // mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_readdatavalid;                                           // mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire  [15:0] mm_interconnect_1_timer_5_s1_writedata;                                  // mm_interconnect_1:timer_5_s1_writedata -> timer_5:writedata
	wire   [2:0] mm_interconnect_1_timer_5_s1_address;                                    // mm_interconnect_1:timer_5_s1_address -> timer_5:address
	wire         mm_interconnect_1_timer_5_s1_chipselect;                                 // mm_interconnect_1:timer_5_s1_chipselect -> timer_5:chipselect
	wire         mm_interconnect_1_timer_5_s1_write;                                      // mm_interconnect_1:timer_5_s1_write -> timer_5:write_n
	wire  [15:0] mm_interconnect_1_timer_5_s1_readdata;                                   // timer_5:readdata -> mm_interconnect_1:timer_5_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_7_s1_writedata;                                  // mm_interconnect_1:timer_7_s1_writedata -> timer_7:writedata
	wire   [2:0] mm_interconnect_1_timer_7_s1_address;                                    // mm_interconnect_1:timer_7_s1_address -> timer_7:address
	wire         mm_interconnect_1_timer_7_s1_chipselect;                                 // mm_interconnect_1:timer_7_s1_chipselect -> timer_7:chipselect
	wire         mm_interconnect_1_timer_7_s1_write;                                      // mm_interconnect_1:timer_7_s1_write -> timer_7:write_n
	wire  [15:0] mm_interconnect_1_timer_7_s1_readdata;                                   // timer_7:readdata -> mm_interconnect_1:timer_7_s1_readdata
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_writedata;                                   // mm_interconnect_1:sd_cmd_s1_writedata -> sd_cmd:writedata
	wire   [1:0] mm_interconnect_1_sd_cmd_s1_address;                                     // mm_interconnect_1:sd_cmd_s1_address -> sd_cmd:address
	wire         mm_interconnect_1_sd_cmd_s1_chipselect;                                  // mm_interconnect_1:sd_cmd_s1_chipselect -> sd_cmd:chipselect
	wire         mm_interconnect_1_sd_cmd_s1_write;                                       // mm_interconnect_1:sd_cmd_s1_write -> sd_cmd:write_n
	wire  [31:0] mm_interconnect_1_sd_cmd_s1_readdata;                                    // sd_cmd:readdata -> mm_interconnect_1:sd_cmd_s1_readdata
	wire  [31:0] mm_interconnect_1_eep_i2c_sda_s1_writedata;                              // mm_interconnect_1:eep_i2c_sda_s1_writedata -> eep_i2c_sda:writedata
	wire   [1:0] mm_interconnect_1_eep_i2c_sda_s1_address;                                // mm_interconnect_1:eep_i2c_sda_s1_address -> eep_i2c_sda:address
	wire         mm_interconnect_1_eep_i2c_sda_s1_chipselect;                             // mm_interconnect_1:eep_i2c_sda_s1_chipselect -> eep_i2c_sda:chipselect
	wire         mm_interconnect_1_eep_i2c_sda_s1_write;                                  // mm_interconnect_1:eep_i2c_sda_s1_write -> eep_i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_eep_i2c_sda_s1_readdata;                               // eep_i2c_sda:readdata -> mm_interconnect_1:eep_i2c_sda_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_8_s1_writedata;                                  // mm_interconnect_1:timer_8_s1_writedata -> timer_8:writedata
	wire   [2:0] mm_interconnect_1_timer_8_s1_address;                                    // mm_interconnect_1:timer_8_s1_address -> timer_8:address
	wire         mm_interconnect_1_timer_8_s1_chipselect;                                 // mm_interconnect_1:timer_8_s1_chipselect -> timer_8:chipselect
	wire         mm_interconnect_1_timer_8_s1_write;                                      // mm_interconnect_1:timer_8_s1_write -> timer_8:write_n
	wire  [15:0] mm_interconnect_1_timer_8_s1_readdata;                                   // timer_8:readdata -> mm_interconnect_1:timer_8_s1_readdata
	wire   [1:0] mm_interconnect_1_ir_s1_address;                                         // mm_interconnect_1:ir_s1_address -> ir:address
	wire  [31:0] mm_interconnect_1_ir_s1_readdata;                                        // ir:readdata -> mm_interconnect_1:ir_s1_readdata
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                                  // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire   [1:0] mm_interconnect_1_i2c_sda_s1_address;                                    // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire         mm_interconnect_1_i2c_sda_s1_chipselect;                                 // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire         mm_interconnect_1_i2c_sda_s1_write;                                      // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire  [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                                   // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;                            // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;                              // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;                           // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire         mm_interconnect_1_sys_clk_timer_s1_write;                                // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;                             // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_writedata;                           // mm_interconnect_1:seg7_avalon_slave_writedata -> seg7:s_writedata
	wire   [2:0] mm_interconnect_1_seg7_avalon_slave_address;                             // mm_interconnect_1:seg7_avalon_slave_address -> seg7:s_address
	wire         mm_interconnect_1_seg7_avalon_slave_write;                               // mm_interconnect_1:seg7_avalon_slave_write -> seg7:s_write
	wire         mm_interconnect_1_seg7_avalon_slave_read;                                // mm_interconnect_1:seg7_avalon_slave_read -> seg7:s_read
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_readdata;                            // seg7:s_readdata -> mm_interconnect_1:seg7_avalon_slave_readdata
	wire  [15:0] mm_interconnect_1_timer_11_s1_writedata;                                 // mm_interconnect_1:timer_11_s1_writedata -> timer_11:writedata
	wire   [2:0] mm_interconnect_1_timer_11_s1_address;                                   // mm_interconnect_1:timer_11_s1_address -> timer_11:address
	wire         mm_interconnect_1_timer_11_s1_chipselect;                                // mm_interconnect_1:timer_11_s1_chipselect -> timer_11:chipselect
	wire         mm_interconnect_1_timer_11_s1_write;                                     // mm_interconnect_1:timer_11_s1_write -> timer_11:write_n
	wire  [15:0] mm_interconnect_1_timer_11_s1_readdata;                                  // timer_11:readdata -> mm_interconnect_1:timer_11_s1_readdata
	wire  [31:0] mm_interconnect_1_ledr_s1_writedata;                                     // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire   [1:0] mm_interconnect_1_ledr_s1_address;                                       // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire         mm_interconnect_1_ledr_s1_chipselect;                                    // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire         mm_interconnect_1_ledr_s1_write;                                         // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_1_ledr_s1_readdata;                                      // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                      // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                        // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_chipselect;                                     // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire         mm_interconnect_1_key_s1_write;                                          // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                       // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_13_s1_writedata;                                 // mm_interconnect_1:timer_13_s1_writedata -> timer_13:writedata
	wire   [2:0] mm_interconnect_1_timer_13_s1_address;                                   // mm_interconnect_1:timer_13_s1_address -> timer_13:address
	wire         mm_interconnect_1_timer_13_s1_chipselect;                                // mm_interconnect_1:timer_13_s1_chipselect -> timer_13:chipselect
	wire         mm_interconnect_1_timer_13_s1_write;                                     // mm_interconnect_1:timer_13_s1_write -> timer_13:write_n
	wire  [15:0] mm_interconnect_1_timer_13_s1_readdata;                                  // timer_13:readdata -> mm_interconnect_1:timer_13_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_10_s1_writedata;                                 // mm_interconnect_1:timer_10_s1_writedata -> timer_10:writedata
	wire   [2:0] mm_interconnect_1_timer_10_s1_address;                                   // mm_interconnect_1:timer_10_s1_address -> timer_10:address
	wire         mm_interconnect_1_timer_10_s1_chipselect;                                // mm_interconnect_1:timer_10_s1_chipselect -> timer_10:chipselect
	wire         mm_interconnect_1_timer_10_s1_write;                                     // mm_interconnect_1:timer_10_s1_write -> timer_10:write_n
	wire  [15:0] mm_interconnect_1_timer_10_s1_readdata;                                  // timer_10:readdata -> mm_interconnect_1:timer_10_s1_readdata
	wire         mm_interconnect_1_sysver_0_avalon_slave_0_waitrequest;                   // sysver_0:waitrequest -> mm_interconnect_1:sysver_0_avalon_slave_0_waitrequest
	wire  [31:0] mm_interconnect_1_sysver_0_avalon_slave_0_writedata;                     // mm_interconnect_1:sysver_0_avalon_slave_0_writedata -> sysver_0:writedata
	wire   [2:0] mm_interconnect_1_sysver_0_avalon_slave_0_address;                       // mm_interconnect_1:sysver_0_avalon_slave_0_address -> sysver_0:address
	wire         mm_interconnect_1_sysver_0_avalon_slave_0_chipselect;                    // mm_interconnect_1:sysver_0_avalon_slave_0_chipselect -> sysver_0:chipselect
	wire         mm_interconnect_1_sysver_0_avalon_slave_0_write;                         // mm_interconnect_1:sysver_0_avalon_slave_0_write -> sysver_0:write
	wire         mm_interconnect_1_sysver_0_avalon_slave_0_read;                          // mm_interconnect_1:sysver_0_avalon_slave_0_read -> sysver_0:read
	wire  [31:0] mm_interconnect_1_sysver_0_avalon_slave_0_readdata;                      // sysver_0:readdata -> mm_interconnect_1:sysver_0_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_1_sysver_0_avalon_slave_0_byteenable;                    // mm_interconnect_1:sysver_0_avalon_slave_0_byteenable -> sysver_0:byteenable
	wire  [15:0] mm_interconnect_1_timer_4_s1_writedata;                                  // mm_interconnect_1:timer_4_s1_writedata -> timer_4:writedata
	wire   [2:0] mm_interconnect_1_timer_4_s1_address;                                    // mm_interconnect_1:timer_4_s1_address -> timer_4:address
	wire         mm_interconnect_1_timer_4_s1_chipselect;                                 // mm_interconnect_1:timer_4_s1_chipselect -> timer_4:chipselect
	wire         mm_interconnect_1_timer_4_s1_write;                                      // mm_interconnect_1:timer_4_s1_write -> timer_4:write_n
	wire  [15:0] mm_interconnect_1_timer_4_s1_readdata;                                   // timer_4:readdata -> mm_interconnect_1:timer_4_s1_readdata
	wire  [31:0] mm_interconnect_1_sd_dat_s1_writedata;                                   // mm_interconnect_1:sd_dat_s1_writedata -> sd_dat:writedata
	wire   [1:0] mm_interconnect_1_sd_dat_s1_address;                                     // mm_interconnect_1:sd_dat_s1_address -> sd_dat:address
	wire         mm_interconnect_1_sd_dat_s1_chipselect;                                  // mm_interconnect_1:sd_dat_s1_chipselect -> sd_dat:chipselect
	wire         mm_interconnect_1_sd_dat_s1_write;                                       // mm_interconnect_1:sd_dat_s1_write -> sd_dat:write_n
	wire  [31:0] mm_interconnect_1_sd_dat_s1_readdata;                                    // sd_dat:readdata -> mm_interconnect_1:sd_dat_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_12_s1_writedata;                                 // mm_interconnect_1:timer_12_s1_writedata -> timer_12:writedata
	wire   [2:0] mm_interconnect_1_timer_12_s1_address;                                   // mm_interconnect_1:timer_12_s1_address -> timer_12:address
	wire         mm_interconnect_1_timer_12_s1_chipselect;                                // mm_interconnect_1:timer_12_s1_chipselect -> timer_12:chipselect
	wire         mm_interconnect_1_timer_12_s1_write;                                     // mm_interconnect_1:timer_12_s1_write -> timer_12:write_n
	wire  [15:0] mm_interconnect_1_timer_12_s1_readdata;                                  // timer_12:readdata -> mm_interconnect_1:timer_12_s1_readdata
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                                  // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire   [1:0] mm_interconnect_1_i2c_scl_s1_address;                                    // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire         mm_interconnect_1_i2c_scl_s1_chipselect;                                 // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire         mm_interconnect_1_i2c_scl_s1_write;                                      // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                                   // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire  [31:0] mm_interconnect_1_eep_i2c_scl_s1_writedata;                              // mm_interconnect_1:eep_i2c_scl_s1_writedata -> eep_i2c_scl:writedata
	wire   [1:0] mm_interconnect_1_eep_i2c_scl_s1_address;                                // mm_interconnect_1:eep_i2c_scl_s1_address -> eep_i2c_scl:address
	wire         mm_interconnect_1_eep_i2c_scl_s1_chipselect;                             // mm_interconnect_1:eep_i2c_scl_s1_chipselect -> eep_i2c_scl:chipselect
	wire         mm_interconnect_1_eep_i2c_scl_s1_write;                                  // mm_interconnect_1:eep_i2c_scl_s1_write -> eep_i2c_scl:write_n
	wire  [31:0] mm_interconnect_1_eep_i2c_scl_s1_readdata;                               // eep_i2c_scl:readdata -> mm_interconnect_1:eep_i2c_scl_s1_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                           // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                          // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire  [15:0] mm_interconnect_1_timer_9_s1_writedata;                                  // mm_interconnect_1:timer_9_s1_writedata -> timer_9:writedata
	wire   [2:0] mm_interconnect_1_timer_9_s1_address;                                    // mm_interconnect_1:timer_9_s1_address -> timer_9:address
	wire         mm_interconnect_1_timer_9_s1_chipselect;                                 // mm_interconnect_1:timer_9_s1_chipselect -> timer_9:chipselect
	wire         mm_interconnect_1_timer_9_s1_write;                                      // mm_interconnect_1:timer_9_s1_write -> timer_9:write_n
	wire  [15:0] mm_interconnect_1_timer_9_s1_readdata;                                   // timer_9:readdata -> mm_interconnect_1:timer_9_s1_readdata
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                                       // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                         // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_chipselect;                                      // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire         mm_interconnect_1_sw_s1_write;                                           // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                        // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [7:0] mm_interconnect_1_lcd_control_slave_writedata;                           // mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	wire   [1:0] mm_interconnect_1_lcd_control_slave_address;                             // mm_interconnect_1:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_1_lcd_control_slave_write;                               // mm_interconnect_1:lcd_control_slave_write -> lcd:write
	wire         mm_interconnect_1_lcd_control_slave_read;                                // mm_interconnect_1:lcd_control_slave_read -> lcd:read
	wire   [7:0] mm_interconnect_1_lcd_control_slave_readdata;                            // lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	wire         mm_interconnect_1_lcd_control_slave_begintransfer;                       // mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire  [15:0] mm_interconnect_1_timer_15_s1_writedata;                                 // mm_interconnect_1:timer_15_s1_writedata -> timer_15:writedata
	wire   [2:0] mm_interconnect_1_timer_15_s1_address;                                   // mm_interconnect_1:timer_15_s1_address -> timer_15:address
	wire         mm_interconnect_1_timer_15_s1_chipselect;                                // mm_interconnect_1:timer_15_s1_chipselect -> timer_15:chipselect
	wire         mm_interconnect_1_timer_15_s1_write;                                     // mm_interconnect_1:timer_15_s1_write -> timer_15:write_n
	wire  [15:0] mm_interconnect_1_timer_15_s1_readdata;                                  // timer_15:readdata -> mm_interconnect_1:timer_15_s1_readdata
	wire  [31:0] mm_interconnect_1_pll_pll_slave_writedata;                               // mm_interconnect_1:pll_pll_slave_writedata -> pll:writedata
	wire   [1:0] mm_interconnect_1_pll_pll_slave_address;                                 // mm_interconnect_1:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_1_pll_pll_slave_write;                                   // mm_interconnect_1:pll_pll_slave_write -> pll:write
	wire         mm_interconnect_1_pll_pll_slave_read;                                    // mm_interconnect_1:pll_pll_slave_read -> pll:read
	wire  [31:0] mm_interconnect_1_pll_pll_slave_readdata;                                // pll:readdata -> mm_interconnect_1:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_1_sd_wp_n_s1_address;                                    // mm_interconnect_1:sd_wp_n_s1_address -> sd_wp_n:address
	wire  [31:0] mm_interconnect_1_sd_wp_n_s1_readdata;                                   // sd_wp_n:readdata -> mm_interconnect_1:sd_wp_n_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_1_s1_writedata;                                  // mm_interconnect_1:timer_1_s1_writedata -> timer_1:writedata
	wire   [2:0] mm_interconnect_1_timer_1_s1_address;                                    // mm_interconnect_1:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_1_timer_1_s1_chipselect;                                 // mm_interconnect_1:timer_1_s1_chipselect -> timer_1:chipselect
	wire         mm_interconnect_1_timer_1_s1_write;                                      // mm_interconnect_1:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_1_timer_1_s1_readdata;                                   // timer_1:readdata -> mm_interconnect_1:timer_1_s1_readdata
	wire  [31:0] mm_interconnect_1_ledg_s1_writedata;                                     // mm_interconnect_1:ledg_s1_writedata -> ledg:writedata
	wire   [1:0] mm_interconnect_1_ledg_s1_address;                                       // mm_interconnect_1:ledg_s1_address -> ledg:address
	wire         mm_interconnect_1_ledg_s1_chipselect;                                    // mm_interconnect_1:ledg_s1_chipselect -> ledg:chipselect
	wire         mm_interconnect_1_ledg_s1_write;                                         // mm_interconnect_1:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_1_ledg_s1_readdata;                                      // ledg:readdata -> mm_interconnect_1:ledg_s1_readdata
	wire  [15:0] mm_interconnect_1_rs232_s1_writedata;                                    // mm_interconnect_1:rs232_s1_writedata -> rs232:writedata
	wire   [2:0] mm_interconnect_1_rs232_s1_address;                                      // mm_interconnect_1:rs232_s1_address -> rs232:address
	wire         mm_interconnect_1_rs232_s1_chipselect;                                   // mm_interconnect_1:rs232_s1_chipselect -> rs232:chipselect
	wire         mm_interconnect_1_rs232_s1_write;                                        // mm_interconnect_1:rs232_s1_write -> rs232:write_n
	wire         mm_interconnect_1_rs232_s1_read;                                         // mm_interconnect_1:rs232_s1_read -> rs232:read_n
	wire  [15:0] mm_interconnect_1_rs232_s1_readdata;                                     // rs232:readdata -> mm_interconnect_1:rs232_s1_readdata
	wire         mm_interconnect_1_rs232_s1_begintransfer;                                // mm_interconnect_1:rs232_s1_begintransfer -> rs232:begintransfer
	wire  [15:0] mm_interconnect_1_timer_6_s1_writedata;                                  // mm_interconnect_1:timer_6_s1_writedata -> timer_6:writedata
	wire   [2:0] mm_interconnect_1_timer_6_s1_address;                                    // mm_interconnect_1:timer_6_s1_address -> timer_6:address
	wire         mm_interconnect_1_timer_6_s1_chipselect;                                 // mm_interconnect_1:timer_6_s1_chipselect -> timer_6:chipselect
	wire         mm_interconnect_1_timer_6_s1_write;                                      // mm_interconnect_1:timer_6_s1_write -> timer_6:write_n
	wire  [15:0] mm_interconnect_1_timer_6_s1_readdata;                                   // timer_6:readdata -> mm_interconnect_1:timer_6_s1_readdata
	wire   [0:0] clock_crossing_io_m0_burstcount;                                         // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire         clock_crossing_io_m0_waitrequest;                                        // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [10:0] clock_crossing_io_m0_address;                                            // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire  [31:0] clock_crossing_io_m0_writedata;                                          // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                              // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire         clock_crossing_io_m0_read;                                               // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire  [31:0] clock_crossing_io_m0_readdata;                                           // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                        // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [3:0] clock_crossing_io_m0_byteenable;                                         // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                      // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [15:0] mm_interconnect_1_timer_0_s1_writedata;                                  // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_1_timer_0_s1_address;                                    // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_1_timer_0_s1_chipselect;                                 // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_1_timer_0_s1_write;                                      // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_1_timer_0_s1_readdata;                                   // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_3_s1_writedata;                                  // mm_interconnect_1:timer_3_s1_writedata -> timer_3:writedata
	wire   [2:0] mm_interconnect_1_timer_3_s1_address;                                    // mm_interconnect_1:timer_3_s1_address -> timer_3:address
	wire         mm_interconnect_1_timer_3_s1_chipselect;                                 // mm_interconnect_1:timer_3_s1_chipselect -> timer_3:chipselect
	wire         mm_interconnect_1_timer_3_s1_write;                                      // mm_interconnect_1:timer_3_s1_write -> timer_3:write_n
	wire  [15:0] mm_interconnect_1_timer_3_s1_readdata;                                   // timer_3:readdata -> mm_interconnect_1:timer_3_s1_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;               // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;                 // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;                // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                      // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                  // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_1_timer_2_s1_writedata;                                  // mm_interconnect_1:timer_2_s1_writedata -> timer_2:writedata
	wire   [2:0] mm_interconnect_1_timer_2_s1_address;                                    // mm_interconnect_1:timer_2_s1_address -> timer_2:address
	wire         mm_interconnect_1_timer_2_s1_chipselect;                                 // mm_interconnect_1:timer_2_s1_chipselect -> timer_2:chipselect
	wire         mm_interconnect_1_timer_2_s1_write;                                      // mm_interconnect_1:timer_2_s1_write -> timer_2:write_n
	wire  [15:0] mm_interconnect_1_timer_2_s1_readdata;                                   // timer_2:readdata -> mm_interconnect_1:timer_2_s1_readdata
	wire  [15:0] mm_interconnect_1_timer_14_s1_writedata;                                 // mm_interconnect_1:timer_14_s1_writedata -> timer_14:writedata
	wire   [2:0] mm_interconnect_1_timer_14_s1_address;                                   // mm_interconnect_1:timer_14_s1_address -> timer_14:address
	wire         mm_interconnect_1_timer_14_s1_chipselect;                                // mm_interconnect_1:timer_14_s1_chipselect -> timer_14:chipselect
	wire         mm_interconnect_1_timer_14_s1_write;                                     // mm_interconnect_1:timer_14_s1_write -> timer_14:write_n
	wire  [15:0] mm_interconnect_1_timer_14_s1_readdata;                                  // timer_14:readdata -> mm_interconnect_1:timer_14_s1_readdata
	wire  [31:0] mm_interconnect_1_sd_clk_s1_writedata;                                   // mm_interconnect_1:sd_clk_s1_writedata -> sd_clk:writedata
	wire   [1:0] mm_interconnect_1_sd_clk_s1_address;                                     // mm_interconnect_1:sd_clk_s1_address -> sd_clk:address
	wire         mm_interconnect_1_sd_clk_s1_chipselect;                                  // mm_interconnect_1:sd_clk_s1_chipselect -> sd_clk:chipselect
	wire         mm_interconnect_1_sd_clk_s1_write;                                       // mm_interconnect_1:sd_clk_s1_write -> sd_clk:write_n
	wire  [31:0] mm_interconnect_1_sd_clk_s1_readdata;                                    // sd_clk:readdata -> mm_interconnect_1:sd_clk_s1_readdata
	wire         irq_mapper_receiver5_irq;                                                // usb:avs_hc_irq_n_oINT0_N -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                // usb:avs_dc_irq_n_oINT0_N -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver24_irq;                                               // uart_0:irq -> irq_mapper:receiver24_irq
	wire         irq_mapper_receiver25_irq;                                               // uart_1:irq -> irq_mapper:receiver25_irq
	wire         irq_mapper_receiver26_irq;                                               // sgdma_rx:csr_irq -> irq_mapper:receiver26_irq
	wire         irq_mapper_receiver27_irq;                                               // sgdma_tx:csr_irq -> irq_mapper:receiver27_irq
	wire  [31:0] vic_0_irq_input_irq;                                                     // irq_mapper:sender_irq -> vic_0:irq_input_irq
	wire         irq_mapper_receiver0_irq;                                                // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                           // sys_clk_timer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                                // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                       // key:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                                // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                       // sw:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                                // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                       // rs232:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver4_irq;                                                // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                       // jtag_uart:av_irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver7_irq;                                                // irq_synchronizer_005:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                                       // timer_0:irq -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver8_irq;                                                // irq_synchronizer_006:sender_irq -> irq_mapper:receiver8_irq
	wire   [0:0] irq_synchronizer_006_receiver_irq;                                       // timer_1:irq -> irq_synchronizer_006:receiver_irq
	wire         irq_mapper_receiver9_irq;                                                // irq_synchronizer_007:sender_irq -> irq_mapper:receiver9_irq
	wire   [0:0] irq_synchronizer_007_receiver_irq;                                       // timer_2:irq -> irq_synchronizer_007:receiver_irq
	wire         irq_mapper_receiver10_irq;                                               // irq_synchronizer_008:sender_irq -> irq_mapper:receiver10_irq
	wire   [0:0] irq_synchronizer_008_receiver_irq;                                       // timer_3:irq -> irq_synchronizer_008:receiver_irq
	wire         irq_mapper_receiver11_irq;                                               // irq_synchronizer_009:sender_irq -> irq_mapper:receiver11_irq
	wire   [0:0] irq_synchronizer_009_receiver_irq;                                       // timer_4:irq -> irq_synchronizer_009:receiver_irq
	wire         irq_mapper_receiver12_irq;                                               // irq_synchronizer_010:sender_irq -> irq_mapper:receiver12_irq
	wire   [0:0] irq_synchronizer_010_receiver_irq;                                       // timer_5:irq -> irq_synchronizer_010:receiver_irq
	wire         irq_mapper_receiver13_irq;                                               // irq_synchronizer_011:sender_irq -> irq_mapper:receiver13_irq
	wire   [0:0] irq_synchronizer_011_receiver_irq;                                       // timer_6:irq -> irq_synchronizer_011:receiver_irq
	wire         irq_mapper_receiver14_irq;                                               // irq_synchronizer_012:sender_irq -> irq_mapper:receiver14_irq
	wire   [0:0] irq_synchronizer_012_receiver_irq;                                       // timer_7:irq -> irq_synchronizer_012:receiver_irq
	wire         irq_mapper_receiver15_irq;                                               // irq_synchronizer_013:sender_irq -> irq_mapper:receiver15_irq
	wire   [0:0] irq_synchronizer_013_receiver_irq;                                       // timer_8:irq -> irq_synchronizer_013:receiver_irq
	wire         irq_mapper_receiver16_irq;                                               // irq_synchronizer_014:sender_irq -> irq_mapper:receiver16_irq
	wire   [0:0] irq_synchronizer_014_receiver_irq;                                       // timer_9:irq -> irq_synchronizer_014:receiver_irq
	wire         irq_mapper_receiver17_irq;                                               // irq_synchronizer_015:sender_irq -> irq_mapper:receiver17_irq
	wire   [0:0] irq_synchronizer_015_receiver_irq;                                       // timer_10:irq -> irq_synchronizer_015:receiver_irq
	wire         irq_mapper_receiver18_irq;                                               // irq_synchronizer_016:sender_irq -> irq_mapper:receiver18_irq
	wire   [0:0] irq_synchronizer_016_receiver_irq;                                       // timer_11:irq -> irq_synchronizer_016:receiver_irq
	wire         irq_mapper_receiver19_irq;                                               // irq_synchronizer_017:sender_irq -> irq_mapper:receiver19_irq
	wire   [0:0] irq_synchronizer_017_receiver_irq;                                       // timer_12:irq -> irq_synchronizer_017:receiver_irq
	wire         irq_mapper_receiver20_irq;                                               // irq_synchronizer_018:sender_irq -> irq_mapper:receiver20_irq
	wire   [0:0] irq_synchronizer_018_receiver_irq;                                       // timer_13:irq -> irq_synchronizer_018:receiver_irq
	wire         irq_mapper_receiver21_irq;                                               // irq_synchronizer_019:sender_irq -> irq_mapper:receiver21_irq
	wire   [0:0] irq_synchronizer_019_receiver_irq;                                       // timer_14:irq -> irq_synchronizer_019:receiver_irq
	wire         irq_mapper_receiver22_irq;                                               // irq_synchronizer_020:sender_irq -> irq_mapper:receiver22_irq
	wire   [0:0] irq_synchronizer_020_receiver_irq;                                       // timer_15:irq -> irq_synchronizer_020:receiver_irq
	wire         irq_mapper_receiver23_irq;                                               // irq_synchronizer_021:sender_irq -> irq_mapper:receiver23_irq
	wire   [0:0] irq_synchronizer_021_receiver_irq;                                       // can_top_0:irq_on -> irq_synchronizer_021:receiver_irq
	wire         tse_receive_endofpacket;                                                 // tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire         tse_receive_valid;                                                       // tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire         tse_receive_startofpacket;                                               // tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire   [5:0] tse_receive_error;                                                       // tse:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_receive_empty;                                                       // tse:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire  [31:0] tse_receive_data;                                                        // tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_receive_ready;                                                       // avalon_st_adapter:in_0_ready -> tse:ff_rx_rdy
	wire         avalon_st_adapter_out_0_endofpacket;                                     // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                           // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire         avalon_st_adapter_out_0_startofpacket;                                   // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                                           // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                                           // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire  [31:0] avalon_st_adapter_out_0_data;                                            // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                                           // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [clock_crossing_io:m0_reset, eep_i2c_scl:reset_n, eep_i2c_sda:reset_n, i2c_scl:reset_n, i2c_sda:reset_n, ir:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, irq_synchronizer_007:receiver_reset, irq_synchronizer_008:receiver_reset, irq_synchronizer_009:receiver_reset, irq_synchronizer_010:receiver_reset, irq_synchronizer_011:receiver_reset, irq_synchronizer_012:receiver_reset, irq_synchronizer_013:receiver_reset, irq_synchronizer_014:receiver_reset, irq_synchronizer_015:receiver_reset, irq_synchronizer_016:receiver_reset, irq_synchronizer_017:receiver_reset, irq_synchronizer_018:receiver_reset, irq_synchronizer_019:receiver_reset, irq_synchronizer_020:receiver_reset, jtag_uart:rst_n, key:reset_n, lcd:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, rs232:reset_n, sd_clk:reset_n, sd_cmd:reset_n, sd_dat:reset_n, sd_wp_n:reset_n, seg7:s_reset, sw:reset_n, sys_clk_timer:reset_n, sysid:reset_n, sysver_0:reset_n, timer_0:reset_n, timer_10:reset_n, timer_11:reset_n, timer_12:reset_n, timer_13:reset_n, timer_14:reset_n, timer_15:reset_n, timer_1:reset_n, timer_2:reset_n, timer_3:reset_n, timer_4:reset_n, timer_5:reset_n, timer_6:reset_n, timer_7:reset_n, timer_8:reset_n, timer_9:reset_n]
	wire         cpu_jtag_debug_module_reset_reset;                                       // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [audio:avs_s1_reset, avalon_st_adapter:in_rst_0_reset, cfi_flash:reset_reset, clock_crossing_io:s0_reset, cpu:reset_n, descriptor_memory:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, irq_synchronizer_008:sender_reset, irq_synchronizer_009:sender_reset, irq_synchronizer_010:sender_reset, irq_synchronizer_011:sender_reset, irq_synchronizer_012:sender_reset, irq_synchronizer_013:sender_reset, irq_synchronizer_014:sender_reset, irq_synchronizer_015:sender_reset, irq_synchronizer_016:sender_reset, irq_synchronizer_017:sender_reset, irq_synchronizer_018:sender_reset, irq_synchronizer_019:sender_reset, irq_synchronizer_020:sender_reset, irq_synchronizer_021:sender_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sdram:reset_n, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sma_in:reset_n, sma_out:reset_n, sram:reset_n, tristate_conduit_bridge_flash:reset, tristate_conduit_pin_sharer_flash:reset_reset, tse:reset, uart_0:reset_n, uart_1:reset_n, usb:avs_dc_reset_n_iRST_N, usb:avs_hc_reset_n_iRST_N, vic_0:clk_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                                  // rst_controller_001:reset_req -> [cpu:reset_req, descriptor_memory:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                      // rst_controller_002:reset_out -> [can_top_0:av_rst_i, irq_synchronizer_021:receiver_reset, mm_interconnect_0:can_top_0_clock_sink_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	DE2_115_SOPC_sys_clk_timer sys_clk_timer (
		.clk        (altpll_io_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                  //   irq.irq
	);

	DE2_115_SOPC_onchip_memory2 onchip_memory2 (
		.clk        (altpll_sys_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	DE2_115_SOPC_sdram sdram (
		.clk            (altpll_sys_clk),                           //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	DE2_115_SOPC_key key (
		.clk        (altpll_io_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)    //                 irq.irq
	);

	DE2_115_SOPC_sma_in sma_in (
		.clk      (altpll_sys_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sma_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sma_in_s1_readdata), //                    .readdata
		.in_port  (sma_in_external_connection_export)     // external_connection.export
	);

	DE2_115_SOPC_sma_out sma_out (
		.clk        (altpll_sys_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_sma_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sma_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sma_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sma_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sma_out_s1_readdata),   //                    .readdata
		.out_port   (sma_out_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sw sw (
		.clk        (altpll_io_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)   //                 irq.irq
	);

	DE2_115_SOPC_ledg ledg (
		.clk        (altpll_io_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_ledr ledr (
		.clk        (altpll_io_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_rs232 rs232 (
		.clk           (altpll_io_clk),                            //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_1_rs232_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_rs232_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_rs232_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_rs232_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_rs232_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_rs232_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_rs232_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (rs232_external_connection_rxd),            // external_connection.export
		.txd           (rs232_external_connection_txd),            //                    .export
		.cts_n         (rs232_external_connection_cts_n),          //                    .export
		.rts_n         (rs232_external_connection_rts_n),          //                    .export
		.irq           (irq_synchronizer_003_receiver_irq)         //                 irq.irq
	);

	DE2_115_SOPC_i2c_scl i2c_scl (
		.clk        (altpll_io_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_i2c_sda i2c_sda (
		.clk        (altpll_io_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_i2c_scl eep_i2c_scl (
		.clk        (altpll_io_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_eep_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_eep_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_eep_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_eep_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_eep_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (eep_i2c_scl_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_i2c_sda eep_i2c_sda (
		.clk        (altpll_io_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_eep_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_eep_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_eep_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_eep_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_eep_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (eep_i2c_sda_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_lcd lcd (
		.reset_n       (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.clk           (altpll_io_clk),                                     //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_control_slave_address),       //              .address
		.LCD_RS        (lcd_external_RS),                                   //      external.export
		.LCD_RW        (lcd_external_RW),                                   //              .export
		.LCD_data      (lcd_external_data),                                 //              .export
		.LCD_E         (lcd_external_E)                                     //              .export
	);

	DE2_115_SOPC_ir ir (
		.clk      (altpll_io_clk),                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_1_ir_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_ir_s1_readdata), //                    .readdata
		.in_port  (ir_external_connection_export)     // external_connection.export
	);

	TERASIC_SRAM #(
		.DATA_BITS (16),
		.ADDR_BITS (20)
	) sram (
		.clk            (altpll_sys_clk),                                  //       clock_reset.clk
		.reset_n        (~rst_controller_001_reset_out_reset),             // clock_reset_reset.reset_n
		.s_chipselect_n (~mm_interconnect_0_sram_avalon_slave_chipselect), //      avalon_slave.chipselect_n
		.s_write_n      (~mm_interconnect_0_sram_avalon_slave_write),      //                  .write_n
		.s_address      (mm_interconnect_0_sram_avalon_slave_address),     //                  .address
		.s_read_n       (~mm_interconnect_0_sram_avalon_slave_read),       //                  .read_n
		.s_writedata    (mm_interconnect_0_sram_avalon_slave_writedata),   //                  .writedata
		.s_readdata     (mm_interconnect_0_sram_avalon_slave_readdata),    //                  .readdata
		.s_byteenable_n (~mm_interconnect_0_sram_avalon_slave_byteenable), //                  .byteenable_n
		.SRAM_DQ        (sram_conduit_end_DQ),                             //       conduit_end.export
		.SRAM_ADDR      (sram_conduit_end_ADDR),                           //                  .export
		.SRAM_UB_n      (sram_conduit_end_UB_n),                           //                  .export
		.SRAM_LB_n      (sram_conduit_end_LB_n),                           //                  .export
		.SRAM_WE_n      (sram_conduit_end_WE_n),                           //                  .export
		.SRAM_CE_n      (sram_conduit_end_CE_n),                           //                  .export
		.SRAM_OE_n      (sram_conduit_end_OE_n)                            //                  .export
	);

	SEG7_IF #(
		.SEG7_NUM       (8),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (mm_interconnect_1_seg7_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_1_seg7_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_1_seg7_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_1_seg7_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_1_seg7_avalon_slave_writedata), //                 .writedata
		.SEG7        (seg7_conduit_end_export),                       //      conduit_end.export
		.s_clk       (altpll_io_clk),                                 //       clock_sink.clk
		.s_reset     (rst_controller_reset_out_reset)                 // clock_sink_reset.reset
	);

	AUDIO_IF audio (
		.avs_s1_address       (mm_interconnect_0_audio_avalon_slave_address),   //     avalon_slave.address
		.avs_s1_read          (mm_interconnect_0_audio_avalon_slave_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_slave_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_0_audio_avalon_slave_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_slave_writedata), //                 .writedata
		.avs_s1_clk           (altpll_sys_clk),                                 //       clock_sink.clk
		.avs_s1_reset         (rst_controller_001_reset_out_reset),             // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                          //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                       //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                       //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                       //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                       //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                          //                 .export
	);

	DE2_115_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_io_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_004_receiver_irq)                          //               irq.irq
	);

	DE2_115_SOPC_i2c_scl sd_clk (
		.clk        (altpll_io_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_sd_clk_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_clk_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_clk_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_clk_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_clk_s1_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_i2c_sda sd_cmd (
		.clk        (altpll_io_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_sd_cmd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_cmd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_cmd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_cmd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_cmd_s1_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_sd_dat sd_dat (
		.clk        (altpll_io_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_1_sd_dat_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_sd_dat_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_sd_dat_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_sd_dat_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_sd_dat_s1_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)       // external_connection.export
	);

	DE2_115_SOPC_ir sd_wp_n (
		.clk      (altpll_io_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_1_sd_wp_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_sd_wp_n_s1_readdata), //                    .readdata
		.in_port  (sd_wp_n_external_connection_export)     // external_connection.export
	);

	DE2_115_SOPC_pll pll (
		.clk       (clk_50_clk),                                //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_1_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_1_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_1_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_1_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_1_pll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_sys_clk),                            //                    c0.clk
		.c1        (altpll_sdram_clk),                          //                    c1.clk
		.c2        (altpll_io_clk),                             //                    c2.clk
		.c3        (altpll_25_clk),                             //                    c3.clk
		.areset    (pll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	ISP1362_IF usb (
		.avs_hc_clk_iCLK           (altpll_sys_clk),                       //       hc_clock.clk
		.avs_hc_reset_n_iRST_N     (~rst_controller_001_reset_out_reset),  // hc_clock_reset.reset_n
		.avs_hc_writedata_iDATA    (mm_interconnect_0_usb_hc_writedata),   //             hc.writedata
		.avs_hc_readdata_oDATA     (mm_interconnect_0_usb_hc_readdata),    //               .readdata
		.avs_hc_address_iADDR      (mm_interconnect_0_usb_hc_address),     //               .address
		.avs_hc_read_n_iRD_N       (~mm_interconnect_0_usb_hc_read),       //               .read_n
		.avs_hc_write_n_iWR_N      (~mm_interconnect_0_usb_hc_write),      //               .write_n
		.avs_hc_chipselect_n_iCS_N (~mm_interconnect_0_usb_hc_chipselect), //               .chipselect_n
		.avs_hc_irq_n_oINT0_N      (irq_mapper_receiver5_irq),             //         hc_irq.irq_n
		.avs_dc_clk_iCLK           (altpll_sys_clk),                       //       dc_clock.clk
		.avs_dc_reset_n_iRST_N     (~rst_controller_001_reset_out_reset),  // dc_clock_reset.reset_n
		.avs_dc_writedata_iDATA    (mm_interconnect_0_usb_dc_writedata),   //             dc.writedata
		.avs_dc_readdata_oDATA     (mm_interconnect_0_usb_dc_readdata),    //               .readdata
		.avs_dc_address_iADDR      (mm_interconnect_0_usb_dc_address),     //               .address
		.avs_dc_read_n_iRD_N       (~mm_interconnect_0_usb_dc_read),       //               .read_n
		.avs_dc_write_n_iWR_N      (~mm_interconnect_0_usb_dc_write),      //               .write_n
		.avs_dc_chipselect_n_iCS_N (~mm_interconnect_0_usb_dc_chipselect), //               .chipselect_n
		.avs_dc_irq_n_oINT0_N      (irq_mapper_receiver6_irq),             //         dc_irq.irq_n
		.USB_DATA                  (usb_conduit_end_DATA),                 //    conduit_end.export
		.USB_ADDR                  (usb_conduit_end_ADDR),                 //               .export
		.USB_RD_N                  (usb_conduit_end_RD_N),                 //               .export
		.USB_WR_N                  (usb_conduit_end_WR_N),                 //               .export
		.USB_CS_N                  (usb_conduit_end_CS_N),                 //               .export
		.USB_RST_N                 (usb_conduit_end_RST_N),                //               .export
		.USB_INT0                  (usb_conduit_end_INT0),                 //               .export
		.USB_INT1                  (usb_conduit_end_INT1)                  //               .export
	);

	sysver #(
		.VER1_ROM_REG_VALUE (32'b00000000000000000000000000000111),
		.VER2_ROM_REG_VALUE (32'b00000000000000000000000000000000),
		.VER3_ROM_REG_VALUE (32'b00000000000000000000000000000001),
		.VER4_ROM_REG_VALUE (32'b00000000000000000000000000000000),
		.VER5_RAM_REG_VALUE (32'b00000000000000000000000000000000),
		.VER6_RAM_REG_VALUE (32'b00000000000000000000000000000000),
		.VER7_RAM_REG_VALUE (32'b00000000000000000000000000000000),
		.VER8_RAM_REG_VALUE (32'b00000000000000000000000000000000)
	) sysver_0 (
		.clk         (altpll_io_clk),                                         //       clock_reset.clk
		.reset_n     (~rst_controller_reset_out_reset),                       // clock_reset_reset.reset_n
		.chipselect  (mm_interconnect_1_sysver_0_avalon_slave_0_chipselect),  //    avalon_slave_0.chipselect
		.address     (mm_interconnect_1_sysver_0_avalon_slave_0_address),     //                  .address
		.write       (mm_interconnect_1_sysver_0_avalon_slave_0_write),       //                  .write
		.writedata   (mm_interconnect_1_sysver_0_avalon_slave_0_writedata),   //                  .writedata
		.read        (mm_interconnect_1_sysver_0_avalon_slave_0_read),        //                  .read
		.readdata    (mm_interconnect_1_sysver_0_avalon_slave_0_readdata),    //                  .readdata
		.byteenable  (mm_interconnect_1_sysver_0_avalon_slave_0_byteenable),  //                  .byteenable
		.waitrequest (mm_interconnect_1_sysver_0_avalon_slave_0_waitrequest)  //                  .waitrequest
	);

	DE2_115_SOPC_sys_clk_timer timer_0 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_005_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_1 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_1_s1_write),     //      .write_n
		.irq        (irq_synchronizer_006_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_2 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_2_s1_write),     //      .write_n
		.irq        (irq_synchronizer_007_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_3 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_3_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_3_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_3_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_3_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_3_s1_write),     //      .write_n
		.irq        (irq_synchronizer_008_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_4 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_4_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_4_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_4_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_4_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_4_s1_write),     //      .write_n
		.irq        (irq_synchronizer_009_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_5 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_5_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_5_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_5_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_5_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_5_s1_write),     //      .write_n
		.irq        (irq_synchronizer_010_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_6 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_6_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_6_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_6_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_6_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_6_s1_write),     //      .write_n
		.irq        (irq_synchronizer_011_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_7 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_7_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_7_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_7_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_7_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_7_s1_write),     //      .write_n
		.irq        (irq_synchronizer_012_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_8 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_8_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_8_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_8_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_8_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_8_s1_write),     //      .write_n
		.irq        (irq_synchronizer_013_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_9 (
		.clk        (altpll_io_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_9_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_9_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_9_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_9_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_9_s1_write),     //      .write_n
		.irq        (irq_synchronizer_014_receiver_irq)        //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_10 (
		.clk        (altpll_io_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_timer_10_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_10_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_10_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_10_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_10_s1_write),     //      .write_n
		.irq        (irq_synchronizer_015_receiver_irq)         //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_11 (
		.clk        (altpll_io_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_timer_11_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_11_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_11_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_11_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_11_s1_write),     //      .write_n
		.irq        (irq_synchronizer_016_receiver_irq)         //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_12 (
		.clk        (altpll_io_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_timer_12_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_12_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_12_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_12_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_12_s1_write),     //      .write_n
		.irq        (irq_synchronizer_017_receiver_irq)         //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_13 (
		.clk        (altpll_io_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_timer_13_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_13_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_13_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_13_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_13_s1_write),     //      .write_n
		.irq        (irq_synchronizer_018_receiver_irq)         //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_14 (
		.clk        (altpll_io_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_timer_14_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_14_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_14_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_14_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_14_s1_write),     //      .write_n
		.irq        (irq_synchronizer_019_receiver_irq)         //   irq.irq
	);

	DE2_115_SOPC_sys_clk_timer timer_15 (
		.clk        (altpll_io_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_timer_15_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_15_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_15_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_15_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_15_s1_write),     //      .write_n
		.irq        (irq_synchronizer_020_receiver_irq)         //   irq.irq
	);

	DE2_115_SOPC_vic_0 vic_0 (
		.clk_clk                        (altpll_sys_clk),                               //                      clk.clk
		.clk_reset_reset                (rst_controller_001_reset_out_reset),           //                clk_reset.reset
		.irq_input_irq                  (vic_0_irq_input_irq),                          //                irq_input.irq
		.csr_access_read                (mm_interconnect_0_vic_0_csr_access_read),      //               csr_access.read
		.csr_access_write               (mm_interconnect_0_vic_0_csr_access_write),     //                         .write
		.csr_access_address             (mm_interconnect_0_vic_0_csr_access_address),   //                         .address
		.csr_access_writedata           (mm_interconnect_0_vic_0_csr_access_writedata), //                         .writedata
		.csr_access_readdata            (mm_interconnect_0_vic_0_csr_access_readdata),  //                         .readdata
		.interrupt_controller_out_valid (vic_0_interrupt_controller_out_valid),         // interrupt_controller_out.valid
		.interrupt_controller_out_data  (vic_0_interrupt_controller_out_data)           //                         .data
	);

	can_top #(
		.Tp (1)
	) can_top_0 (
		.av_cs_i    (mm_interconnect_0_can_top_0_avalon_slave_0_chipselect), //   avalon_slave_0.chipselect
		.av_wr_i    (mm_interconnect_0_can_top_0_avalon_slave_0_write),      //                 .write
		.av_adr_i   (mm_interconnect_0_can_top_0_avalon_slave_0_address),    //                 .address
		.av_dat_i   (mm_interconnect_0_can_top_0_avalon_slave_0_writedata),  //                 .writedata
		.av_dat_o   (mm_interconnect_0_can_top_0_avalon_slave_0_readdata),   //                 .readdata
		.tx_o       (can_top_0_conduit_end_tx_o),                            //      conduit_end.export
		.rx_i       (can_top_0_conduit_end_rx_i),                            //                 .export
		.clkout_o   (can_top_0_conduit_end_clkout_o),                        //                 .export
		.bus_off_on (can_top_0_conduit_end_bus_off_on),                      //                 .export
		.clk_i      (clk_50_clk),                                            //       clock_sink.clk
		.av_rst_i   (rst_controller_002_reset_out_reset),                    // clock_sink_reset.reset
		.irq_on     (irq_synchronizer_021_receiver_irq)                      // interrupt_sender.irq_n
	);

	DE2_115_SOPC_uart_0 uart_0 (
		.clk           (altpll_sys_clk),                            //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver24_irq)                  //                 irq.irq
	);

	DE2_115_SOPC_uart_0 uart_1 (
		.clk           (altpll_sys_clk),                            //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address       (mm_interconnect_0_uart_1_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_1_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_1_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_1_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_1_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_1_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_1_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_1_external_connection_rxd),            // external_connection.export
		.txd           (uart_1_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver25_irq)                  //                 irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (11),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_io_clk),                                        //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (altpll_sys_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SOPC_cpu cpu (
		.clk                                   (altpll_sys_clk),                                      //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_burstcount                          (cpu_instruction_master_burstcount),                   //                          .burstcount
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.eic_port_valid                        (vic_0_interrupt_controller_out_valid),                //   interrupt_controller_in.valid
		.eic_port_data                         (vic_0_interrupt_controller_out_data),                 //                          .data
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE2_115_SOPC_sysid sysid (
		.clock    (altpll_io_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE2_115_SOPC_tristate_conduit_bridge_flash tristate_conduit_bridge_flash (
		.clk                                   (altpll_sys_clk),                                                          //   clk.clk
		.reset                                 (rst_controller_001_reset_out_reset),                                      // reset.reset
		.request                               (tristate_conduit_pin_sharer_flash_tcm_request),                           //   tcs.request
		.grant                                 (tristate_conduit_pin_sharer_flash_tcm_grant),                             //      .grant
		.tcs_address_to_the_cfi_flash          (tristate_conduit_pin_sharer_flash_tcm_address_to_the_cfi_flash_out),      //      .address_to_the_cfi_flash_out
		.tcs_tri_state_bridge_flash_data       (tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_out),   //      .tri_state_bridge_flash_data_out
		.tcs_tri_state_bridge_flash_data_outen (tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_outen), //      .tri_state_bridge_flash_data_outen
		.tcs_tri_state_bridge_flash_data_in    (tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_in),    //      .tri_state_bridge_flash_data_in
		.tcs_write_n_to_the_cfi_flash          (tristate_conduit_pin_sharer_flash_tcm_write_n_to_the_cfi_flash_out),      //      .write_n_to_the_cfi_flash_out
		.tcs_select_n_to_the_cfi_flash         (tristate_conduit_pin_sharer_flash_tcm_select_n_to_the_cfi_flash_out),     //      .select_n_to_the_cfi_flash_out
		.tcs_read_n_to_the_cfi_flash           (tristate_conduit_pin_sharer_flash_tcm_read_n_to_the_cfi_flash_out),       //      .read_n_to_the_cfi_flash_out
		.address_to_the_cfi_flash              (tristate_conduit_bridge_flash_out_address_to_the_cfi_flash),              //   out.address_to_the_cfi_flash
		.tri_state_bridge_flash_data           (tristate_conduit_bridge_flash_out_tri_state_bridge_flash_data),           //      .tri_state_bridge_flash_data
		.write_n_to_the_cfi_flash              (tristate_conduit_bridge_flash_out_write_n_to_the_cfi_flash),              //      .write_n_to_the_cfi_flash
		.select_n_to_the_cfi_flash             (tristate_conduit_bridge_flash_out_select_n_to_the_cfi_flash),             //      .select_n_to_the_cfi_flash
		.read_n_to_the_cfi_flash               (tristate_conduit_bridge_flash_out_read_n_to_the_cfi_flash)                //      .read_n_to_the_cfi_flash
	);

	DE2_115_SOPC_tristate_conduit_pin_sharer_flash tristate_conduit_pin_sharer_flash (
		.clk_clk                           (altpll_sys_clk),                                                          //   clk.clk
		.reset_reset                       (rst_controller_001_reset_out_reset),                                      // reset.reset
		.request                           (tristate_conduit_pin_sharer_flash_tcm_request),                           //   tcm.request
		.grant                             (tristate_conduit_pin_sharer_flash_tcm_grant),                             //      .grant
		.address_to_the_cfi_flash          (tristate_conduit_pin_sharer_flash_tcm_address_to_the_cfi_flash_out),      //      .address_to_the_cfi_flash_out
		.read_n_to_the_cfi_flash           (tristate_conduit_pin_sharer_flash_tcm_read_n_to_the_cfi_flash_out),       //      .read_n_to_the_cfi_flash_out
		.write_n_to_the_cfi_flash          (tristate_conduit_pin_sharer_flash_tcm_write_n_to_the_cfi_flash_out),      //      .write_n_to_the_cfi_flash_out
		.tri_state_bridge_flash_data       (tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_out),   //      .tri_state_bridge_flash_data_out
		.tri_state_bridge_flash_data_in    (tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_in),    //      .tri_state_bridge_flash_data_in
		.tri_state_bridge_flash_data_outen (tristate_conduit_pin_sharer_flash_tcm_tri_state_bridge_flash_data_outen), //      .tri_state_bridge_flash_data_outen
		.select_n_to_the_cfi_flash         (tristate_conduit_pin_sharer_flash_tcm_select_n_to_the_cfi_flash_out),     //      .select_n_to_the_cfi_flash_out
		.tcs0_request                      (cfi_flash_tcm_request),                                                   //  tcs0.request
		.tcs0_grant                        (cfi_flash_tcm_grant),                                                     //      .grant
		.tcs0_address_out                  (cfi_flash_tcm_address_out),                                               //      .address_out
		.tcs0_read_n_out                   (cfi_flash_tcm_read_n_out),                                                //      .read_n_out
		.tcs0_write_n_out                  (cfi_flash_tcm_write_n_out),                                               //      .write_n_out
		.tcs0_data_out                     (cfi_flash_tcm_data_out),                                                  //      .data_out
		.tcs0_data_in                      (cfi_flash_tcm_data_in),                                                   //      .data_in
		.tcs0_data_outen                   (cfi_flash_tcm_data_outen),                                                //      .data_outen
		.tcs0_chipselect_n_out             (cfi_flash_tcm_chipselect_n_out)                                           //      .chipselect_n_out
	);

	DE2_115_SOPC_cfi_flash #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash (
		.clk_clk              (altpll_sys_clk),                                //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),            // reset.reset
		.uas_address          (mm_interconnect_0_cfi_flash_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_cfi_flash_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_cfi_flash_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_cfi_flash_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_cfi_flash_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_cfi_flash_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_cfi_flash_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_cfi_flash_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_cfi_flash_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_cfi_flash_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_cfi_flash_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (cfi_flash_tcm_request),                         //      .request
		.tcm_grant            (cfi_flash_tcm_grant),                           //      .grant
		.tcm_address_out      (cfi_flash_tcm_address_out),                     //      .address_out
		.tcm_data_out         (cfi_flash_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (cfi_flash_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (cfi_flash_tcm_data_in)                          //      .data_in
	);

	DE2_115_SOPC_tse tse (
		.clk           (altpll_sys_clk),                                 // control_port_clock_connection.clk
		.reset         (rst_controller_001_reset_out_reset),             //              reset_connection.reset
		.address       (mm_interconnect_0_tse_control_port_address),     //                  control_port.address
		.readdata      (mm_interconnect_0_tse_control_port_readdata),    //                              .readdata
		.read          (mm_interconnect_0_tse_control_port_read),        //                              .read
		.writedata     (mm_interconnect_0_tse_control_port_writedata),   //                              .writedata
		.write         (mm_interconnect_0_tse_control_port_write),       //                              .write
		.waitrequest   (mm_interconnect_0_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (tse_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (tse_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (tse_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (tse_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (tse_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (tse_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (tse_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (altpll_sys_clk),                                 //      receive_clock_connection.clk
		.ff_tx_clk     (altpll_sys_clk),                                 //     transmit_clock_connection.clk
		.ff_rx_data    (tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_receive_error),                              //                              .error
		.ff_rx_mod     (tse_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                              //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                       //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                             //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                             //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                             //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                     //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                             //                              .valid
		.mdc           (tse_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (tse_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (tse_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (tse_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.ff_tx_crc_fwd (tse_mac_misc_connection_ff_tx_crc_fwd),          //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy   (tse_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (tse_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (tse_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (tse_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (tse_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (tse_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (tse_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (tse_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (tse_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	DE2_115_SOPC_sgdma_rx sgdma_rx (
		.clk                           (altpll_sys_clk),                            //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver26_irq),                 //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	DE2_115_SOPC_sgdma_tx sgdma_tx (
		.clk                           (altpll_sys_clk),                            //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver27_irq),                 //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	DE2_115_SOPC_descriptor_memory descriptor_memory (
		.clk        (altpll_sys_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)             //       .reset_req
	);

	DE2_115_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                         (clk_50_clk),                                            //                                       clk_50_clk.clk
		.pll_c0_clk                                             (altpll_sys_clk),                                        //                                           pll_c0.clk
		.can_top_0_clock_sink_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                    // can_top_0_clock_sink_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                    //                cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                                (cpu_data_master_address),                               //                                  cpu_data_master.address
		.cpu_data_master_waitrequest                            (cpu_data_master_waitrequest),                           //                                                 .waitrequest
		.cpu_data_master_byteenable                             (cpu_data_master_byteenable),                            //                                                 .byteenable
		.cpu_data_master_read                                   (cpu_data_master_read),                                  //                                                 .read
		.cpu_data_master_readdata                               (cpu_data_master_readdata),                              //                                                 .readdata
		.cpu_data_master_write                                  (cpu_data_master_write),                                 //                                                 .write
		.cpu_data_master_writedata                              (cpu_data_master_writedata),                             //                                                 .writedata
		.cpu_data_master_debugaccess                            (cpu_data_master_debugaccess),                           //                                                 .debugaccess
		.cpu_instruction_master_address                         (cpu_instruction_master_address),                        //                           cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                     (cpu_instruction_master_waitrequest),                    //                                                 .waitrequest
		.cpu_instruction_master_burstcount                      (cpu_instruction_master_burstcount),                     //                                                 .burstcount
		.cpu_instruction_master_read                            (cpu_instruction_master_read),                           //                                                 .read
		.cpu_instruction_master_readdata                        (cpu_instruction_master_readdata),                       //                                                 .readdata
		.cpu_instruction_master_readdatavalid                   (cpu_instruction_master_readdatavalid),                  //                                                 .readdatavalid
		.sgdma_rx_descriptor_read_address                       (sgdma_rx_descriptor_read_address),                      //                         sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest                   (sgdma_rx_descriptor_read_waitrequest),                  //                                                 .waitrequest
		.sgdma_rx_descriptor_read_read                          (sgdma_rx_descriptor_read_read),                         //                                                 .read
		.sgdma_rx_descriptor_read_readdata                      (sgdma_rx_descriptor_read_readdata),                     //                                                 .readdata
		.sgdma_rx_descriptor_read_readdatavalid                 (sgdma_rx_descriptor_read_readdatavalid),                //                                                 .readdatavalid
		.sgdma_rx_descriptor_write_address                      (sgdma_rx_descriptor_write_address),                     //                        sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest                  (sgdma_rx_descriptor_write_waitrequest),                 //                                                 .waitrequest
		.sgdma_rx_descriptor_write_write                        (sgdma_rx_descriptor_write_write),                       //                                                 .write
		.sgdma_rx_descriptor_write_writedata                    (sgdma_rx_descriptor_write_writedata),                   //                                                 .writedata
		.sgdma_rx_m_write_address                               (sgdma_rx_m_write_address),                              //                                 sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest                           (sgdma_rx_m_write_waitrequest),                          //                                                 .waitrequest
		.sgdma_rx_m_write_byteenable                            (sgdma_rx_m_write_byteenable),                           //                                                 .byteenable
		.sgdma_rx_m_write_write                                 (sgdma_rx_m_write_write),                                //                                                 .write
		.sgdma_rx_m_write_writedata                             (sgdma_rx_m_write_writedata),                            //                                                 .writedata
		.sgdma_tx_descriptor_read_address                       (sgdma_tx_descriptor_read_address),                      //                         sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest                   (sgdma_tx_descriptor_read_waitrequest),                  //                                                 .waitrequest
		.sgdma_tx_descriptor_read_read                          (sgdma_tx_descriptor_read_read),                         //                                                 .read
		.sgdma_tx_descriptor_read_readdata                      (sgdma_tx_descriptor_read_readdata),                     //                                                 .readdata
		.sgdma_tx_descriptor_read_readdatavalid                 (sgdma_tx_descriptor_read_readdatavalid),                //                                                 .readdatavalid
		.sgdma_tx_descriptor_write_address                      (sgdma_tx_descriptor_write_address),                     //                        sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest                  (sgdma_tx_descriptor_write_waitrequest),                 //                                                 .waitrequest
		.sgdma_tx_descriptor_write_write                        (sgdma_tx_descriptor_write_write),                       //                                                 .write
		.sgdma_tx_descriptor_write_writedata                    (sgdma_tx_descriptor_write_writedata),                   //                                                 .writedata
		.sgdma_tx_m_read_address                                (sgdma_tx_m_read_address),                               //                                  sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest                            (sgdma_tx_m_read_waitrequest),                           //                                                 .waitrequest
		.sgdma_tx_m_read_read                                   (sgdma_tx_m_read_read),                                  //                                                 .read
		.sgdma_tx_m_read_readdata                               (sgdma_tx_m_read_readdata),                              //                                                 .readdata
		.sgdma_tx_m_read_readdatavalid                          (sgdma_tx_m_read_readdatavalid),                         //                                                 .readdatavalid
		.audio_avalon_slave_address                             (mm_interconnect_0_audio_avalon_slave_address),          //                               audio_avalon_slave.address
		.audio_avalon_slave_write                               (mm_interconnect_0_audio_avalon_slave_write),            //                                                 .write
		.audio_avalon_slave_read                                (mm_interconnect_0_audio_avalon_slave_read),             //                                                 .read
		.audio_avalon_slave_readdata                            (mm_interconnect_0_audio_avalon_slave_readdata),         //                                                 .readdata
		.audio_avalon_slave_writedata                           (mm_interconnect_0_audio_avalon_slave_writedata),        //                                                 .writedata
		.can_top_0_avalon_slave_0_address                       (mm_interconnect_0_can_top_0_avalon_slave_0_address),    //                         can_top_0_avalon_slave_0.address
		.can_top_0_avalon_slave_0_write                         (mm_interconnect_0_can_top_0_avalon_slave_0_write),      //                                                 .write
		.can_top_0_avalon_slave_0_readdata                      (mm_interconnect_0_can_top_0_avalon_slave_0_readdata),   //                                                 .readdata
		.can_top_0_avalon_slave_0_writedata                     (mm_interconnect_0_can_top_0_avalon_slave_0_writedata),  //                                                 .writedata
		.can_top_0_avalon_slave_0_chipselect                    (mm_interconnect_0_can_top_0_avalon_slave_0_chipselect), //                                                 .chipselect
		.cfi_flash_uas_address                                  (mm_interconnect_0_cfi_flash_uas_address),               //                                    cfi_flash_uas.address
		.cfi_flash_uas_write                                    (mm_interconnect_0_cfi_flash_uas_write),                 //                                                 .write
		.cfi_flash_uas_read                                     (mm_interconnect_0_cfi_flash_uas_read),                  //                                                 .read
		.cfi_flash_uas_readdata                                 (mm_interconnect_0_cfi_flash_uas_readdata),              //                                                 .readdata
		.cfi_flash_uas_writedata                                (mm_interconnect_0_cfi_flash_uas_writedata),             //                                                 .writedata
		.cfi_flash_uas_burstcount                               (mm_interconnect_0_cfi_flash_uas_burstcount),            //                                                 .burstcount
		.cfi_flash_uas_byteenable                               (mm_interconnect_0_cfi_flash_uas_byteenable),            //                                                 .byteenable
		.cfi_flash_uas_readdatavalid                            (mm_interconnect_0_cfi_flash_uas_readdatavalid),         //                                                 .readdatavalid
		.cfi_flash_uas_waitrequest                              (mm_interconnect_0_cfi_flash_uas_waitrequest),           //                                                 .waitrequest
		.cfi_flash_uas_lock                                     (mm_interconnect_0_cfi_flash_uas_lock),                  //                                                 .lock
		.cfi_flash_uas_debugaccess                              (mm_interconnect_0_cfi_flash_uas_debugaccess),           //                                                 .debugaccess
		.clock_crossing_io_s0_address                           (mm_interconnect_0_clock_crossing_io_s0_address),        //                             clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                             (mm_interconnect_0_clock_crossing_io_s0_write),          //                                                 .write
		.clock_crossing_io_s0_read                              (mm_interconnect_0_clock_crossing_io_s0_read),           //                                                 .read
		.clock_crossing_io_s0_readdata                          (mm_interconnect_0_clock_crossing_io_s0_readdata),       //                                                 .readdata
		.clock_crossing_io_s0_writedata                         (mm_interconnect_0_clock_crossing_io_s0_writedata),      //                                                 .writedata
		.clock_crossing_io_s0_burstcount                        (mm_interconnect_0_clock_crossing_io_s0_burstcount),     //                                                 .burstcount
		.clock_crossing_io_s0_byteenable                        (mm_interconnect_0_clock_crossing_io_s0_byteenable),     //                                                 .byteenable
		.clock_crossing_io_s0_readdatavalid                     (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),  //                                                 .readdatavalid
		.clock_crossing_io_s0_waitrequest                       (mm_interconnect_0_clock_crossing_io_s0_waitrequest),    //                                                 .waitrequest
		.clock_crossing_io_s0_debugaccess                       (mm_interconnect_0_clock_crossing_io_s0_debugaccess),    //                                                 .debugaccess
		.cpu_jtag_debug_module_address                          (mm_interconnect_0_cpu_jtag_debug_module_address),       //                            cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                            (mm_interconnect_0_cpu_jtag_debug_module_write),         //                                                 .write
		.cpu_jtag_debug_module_read                             (mm_interconnect_0_cpu_jtag_debug_module_read),          //                                                 .read
		.cpu_jtag_debug_module_readdata                         (mm_interconnect_0_cpu_jtag_debug_module_readdata),      //                                                 .readdata
		.cpu_jtag_debug_module_writedata                        (mm_interconnect_0_cpu_jtag_debug_module_writedata),     //                                                 .writedata
		.cpu_jtag_debug_module_byteenable                       (mm_interconnect_0_cpu_jtag_debug_module_byteenable),    //                                                 .byteenable
		.cpu_jtag_debug_module_waitrequest                      (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),   //                                                 .waitrequest
		.cpu_jtag_debug_module_debugaccess                      (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),   //                                                 .debugaccess
		.descriptor_memory_s1_address                           (mm_interconnect_0_descriptor_memory_s1_address),        //                             descriptor_memory_s1.address
		.descriptor_memory_s1_write                             (mm_interconnect_0_descriptor_memory_s1_write),          //                                                 .write
		.descriptor_memory_s1_readdata                          (mm_interconnect_0_descriptor_memory_s1_readdata),       //                                                 .readdata
		.descriptor_memory_s1_writedata                         (mm_interconnect_0_descriptor_memory_s1_writedata),      //                                                 .writedata
		.descriptor_memory_s1_byteenable                        (mm_interconnect_0_descriptor_memory_s1_byteenable),     //                                                 .byteenable
		.descriptor_memory_s1_chipselect                        (mm_interconnect_0_descriptor_memory_s1_chipselect),     //                                                 .chipselect
		.descriptor_memory_s1_clken                             (mm_interconnect_0_descriptor_memory_s1_clken),          //                                                 .clken
		.onchip_memory2_s1_address                              (mm_interconnect_0_onchip_memory2_s1_address),           //                                onchip_memory2_s1.address
		.onchip_memory2_s1_write                                (mm_interconnect_0_onchip_memory2_s1_write),             //                                                 .write
		.onchip_memory2_s1_readdata                             (mm_interconnect_0_onchip_memory2_s1_readdata),          //                                                 .readdata
		.onchip_memory2_s1_writedata                            (mm_interconnect_0_onchip_memory2_s1_writedata),         //                                                 .writedata
		.onchip_memory2_s1_byteenable                           (mm_interconnect_0_onchip_memory2_s1_byteenable),        //                                                 .byteenable
		.onchip_memory2_s1_chipselect                           (mm_interconnect_0_onchip_memory2_s1_chipselect),        //                                                 .chipselect
		.onchip_memory2_s1_clken                                (mm_interconnect_0_onchip_memory2_s1_clken),             //                                                 .clken
		.sdram_s1_address                                       (mm_interconnect_0_sdram_s1_address),                    //                                         sdram_s1.address
		.sdram_s1_write                                         (mm_interconnect_0_sdram_s1_write),                      //                                                 .write
		.sdram_s1_read                                          (mm_interconnect_0_sdram_s1_read),                       //                                                 .read
		.sdram_s1_readdata                                      (mm_interconnect_0_sdram_s1_readdata),                   //                                                 .readdata
		.sdram_s1_writedata                                     (mm_interconnect_0_sdram_s1_writedata),                  //                                                 .writedata
		.sdram_s1_byteenable                                    (mm_interconnect_0_sdram_s1_byteenable),                 //                                                 .byteenable
		.sdram_s1_readdatavalid                                 (mm_interconnect_0_sdram_s1_readdatavalid),              //                                                 .readdatavalid
		.sdram_s1_waitrequest                                   (mm_interconnect_0_sdram_s1_waitrequest),                //                                                 .waitrequest
		.sdram_s1_chipselect                                    (mm_interconnect_0_sdram_s1_chipselect),                 //                                                 .chipselect
		.sgdma_rx_csr_address                                   (mm_interconnect_0_sgdma_rx_csr_address),                //                                     sgdma_rx_csr.address
		.sgdma_rx_csr_write                                     (mm_interconnect_0_sgdma_rx_csr_write),                  //                                                 .write
		.sgdma_rx_csr_read                                      (mm_interconnect_0_sgdma_rx_csr_read),                   //                                                 .read
		.sgdma_rx_csr_readdata                                  (mm_interconnect_0_sgdma_rx_csr_readdata),               //                                                 .readdata
		.sgdma_rx_csr_writedata                                 (mm_interconnect_0_sgdma_rx_csr_writedata),              //                                                 .writedata
		.sgdma_rx_csr_chipselect                                (mm_interconnect_0_sgdma_rx_csr_chipselect),             //                                                 .chipselect
		.sgdma_tx_csr_address                                   (mm_interconnect_0_sgdma_tx_csr_address),                //                                     sgdma_tx_csr.address
		.sgdma_tx_csr_write                                     (mm_interconnect_0_sgdma_tx_csr_write),                  //                                                 .write
		.sgdma_tx_csr_read                                      (mm_interconnect_0_sgdma_tx_csr_read),                   //                                                 .read
		.sgdma_tx_csr_readdata                                  (mm_interconnect_0_sgdma_tx_csr_readdata),               //                                                 .readdata
		.sgdma_tx_csr_writedata                                 (mm_interconnect_0_sgdma_tx_csr_writedata),              //                                                 .writedata
		.sgdma_tx_csr_chipselect                                (mm_interconnect_0_sgdma_tx_csr_chipselect),             //                                                 .chipselect
		.sma_in_s1_address                                      (mm_interconnect_0_sma_in_s1_address),                   //                                        sma_in_s1.address
		.sma_in_s1_readdata                                     (mm_interconnect_0_sma_in_s1_readdata),                  //                                                 .readdata
		.sma_out_s1_address                                     (mm_interconnect_0_sma_out_s1_address),                  //                                       sma_out_s1.address
		.sma_out_s1_write                                       (mm_interconnect_0_sma_out_s1_write),                    //                                                 .write
		.sma_out_s1_readdata                                    (mm_interconnect_0_sma_out_s1_readdata),                 //                                                 .readdata
		.sma_out_s1_writedata                                   (mm_interconnect_0_sma_out_s1_writedata),                //                                                 .writedata
		.sma_out_s1_chipselect                                  (mm_interconnect_0_sma_out_s1_chipselect),               //                                                 .chipselect
		.sram_avalon_slave_address                              (mm_interconnect_0_sram_avalon_slave_address),           //                                sram_avalon_slave.address
		.sram_avalon_slave_write                                (mm_interconnect_0_sram_avalon_slave_write),             //                                                 .write
		.sram_avalon_slave_read                                 (mm_interconnect_0_sram_avalon_slave_read),              //                                                 .read
		.sram_avalon_slave_readdata                             (mm_interconnect_0_sram_avalon_slave_readdata),          //                                                 .readdata
		.sram_avalon_slave_writedata                            (mm_interconnect_0_sram_avalon_slave_writedata),         //                                                 .writedata
		.sram_avalon_slave_byteenable                           (mm_interconnect_0_sram_avalon_slave_byteenable),        //                                                 .byteenable
		.sram_avalon_slave_chipselect                           (mm_interconnect_0_sram_avalon_slave_chipselect),        //                                                 .chipselect
		.tse_control_port_address                               (mm_interconnect_0_tse_control_port_address),            //                                 tse_control_port.address
		.tse_control_port_write                                 (mm_interconnect_0_tse_control_port_write),              //                                                 .write
		.tse_control_port_read                                  (mm_interconnect_0_tse_control_port_read),               //                                                 .read
		.tse_control_port_readdata                              (mm_interconnect_0_tse_control_port_readdata),           //                                                 .readdata
		.tse_control_port_writedata                             (mm_interconnect_0_tse_control_port_writedata),          //                                                 .writedata
		.tse_control_port_waitrequest                           (mm_interconnect_0_tse_control_port_waitrequest),        //                                                 .waitrequest
		.uart_0_s1_address                                      (mm_interconnect_0_uart_0_s1_address),                   //                                        uart_0_s1.address
		.uart_0_s1_write                                        (mm_interconnect_0_uart_0_s1_write),                     //                                                 .write
		.uart_0_s1_read                                         (mm_interconnect_0_uart_0_s1_read),                      //                                                 .read
		.uart_0_s1_readdata                                     (mm_interconnect_0_uart_0_s1_readdata),                  //                                                 .readdata
		.uart_0_s1_writedata                                    (mm_interconnect_0_uart_0_s1_writedata),                 //                                                 .writedata
		.uart_0_s1_begintransfer                                (mm_interconnect_0_uart_0_s1_begintransfer),             //                                                 .begintransfer
		.uart_0_s1_chipselect                                   (mm_interconnect_0_uart_0_s1_chipselect),                //                                                 .chipselect
		.uart_1_s1_address                                      (mm_interconnect_0_uart_1_s1_address),                   //                                        uart_1_s1.address
		.uart_1_s1_write                                        (mm_interconnect_0_uart_1_s1_write),                     //                                                 .write
		.uart_1_s1_read                                         (mm_interconnect_0_uart_1_s1_read),                      //                                                 .read
		.uart_1_s1_readdata                                     (mm_interconnect_0_uart_1_s1_readdata),                  //                                                 .readdata
		.uart_1_s1_writedata                                    (mm_interconnect_0_uart_1_s1_writedata),                 //                                                 .writedata
		.uart_1_s1_begintransfer                                (mm_interconnect_0_uart_1_s1_begintransfer),             //                                                 .begintransfer
		.uart_1_s1_chipselect                                   (mm_interconnect_0_uart_1_s1_chipselect),                //                                                 .chipselect
		.usb_dc_address                                         (mm_interconnect_0_usb_dc_address),                      //                                           usb_dc.address
		.usb_dc_write                                           (mm_interconnect_0_usb_dc_write),                        //                                                 .write
		.usb_dc_read                                            (mm_interconnect_0_usb_dc_read),                         //                                                 .read
		.usb_dc_readdata                                        (mm_interconnect_0_usb_dc_readdata),                     //                                                 .readdata
		.usb_dc_writedata                                       (mm_interconnect_0_usb_dc_writedata),                    //                                                 .writedata
		.usb_dc_chipselect                                      (mm_interconnect_0_usb_dc_chipselect),                   //                                                 .chipselect
		.usb_hc_address                                         (mm_interconnect_0_usb_hc_address),                      //                                           usb_hc.address
		.usb_hc_write                                           (mm_interconnect_0_usb_hc_write),                        //                                                 .write
		.usb_hc_read                                            (mm_interconnect_0_usb_hc_read),                         //                                                 .read
		.usb_hc_readdata                                        (mm_interconnect_0_usb_hc_readdata),                     //                                                 .readdata
		.usb_hc_writedata                                       (mm_interconnect_0_usb_hc_writedata),                    //                                                 .writedata
		.usb_hc_chipselect                                      (mm_interconnect_0_usb_hc_chipselect),                   //                                                 .chipselect
		.vic_0_csr_access_address                               (mm_interconnect_0_vic_0_csr_access_address),            //                                 vic_0_csr_access.address
		.vic_0_csr_access_write                                 (mm_interconnect_0_vic_0_csr_access_write),              //                                                 .write
		.vic_0_csr_access_read                                  (mm_interconnect_0_vic_0_csr_access_read),               //                                                 .read
		.vic_0_csr_access_readdata                              (mm_interconnect_0_vic_0_csr_access_readdata),           //                                                 .readdata
		.vic_0_csr_access_writedata                             (mm_interconnect_0_vic_0_csr_access_writedata)           //                                                 .writedata
	);

	DE2_115_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.clk_50_clk_clk                                         (clk_50_clk),                                                //                                       clk_50_clk.clk
		.pll_c2_clk                                             (altpll_io_clk),                                             //                                           pll_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset  (rst_controller_002_reset_out_reset),                        //  pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                              //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                          //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                           //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                           //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                                 //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                             //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),                        //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                                //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                            //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                          //                                                 .debugaccess
		.eep_i2c_scl_s1_address                                 (mm_interconnect_1_eep_i2c_scl_s1_address),                  //                                   eep_i2c_scl_s1.address
		.eep_i2c_scl_s1_write                                   (mm_interconnect_1_eep_i2c_scl_s1_write),                    //                                                 .write
		.eep_i2c_scl_s1_readdata                                (mm_interconnect_1_eep_i2c_scl_s1_readdata),                 //                                                 .readdata
		.eep_i2c_scl_s1_writedata                               (mm_interconnect_1_eep_i2c_scl_s1_writedata),                //                                                 .writedata
		.eep_i2c_scl_s1_chipselect                              (mm_interconnect_1_eep_i2c_scl_s1_chipselect),               //                                                 .chipselect
		.eep_i2c_sda_s1_address                                 (mm_interconnect_1_eep_i2c_sda_s1_address),                  //                                   eep_i2c_sda_s1.address
		.eep_i2c_sda_s1_write                                   (mm_interconnect_1_eep_i2c_sda_s1_write),                    //                                                 .write
		.eep_i2c_sda_s1_readdata                                (mm_interconnect_1_eep_i2c_sda_s1_readdata),                 //                                                 .readdata
		.eep_i2c_sda_s1_writedata                               (mm_interconnect_1_eep_i2c_sda_s1_writedata),                //                                                 .writedata
		.eep_i2c_sda_s1_chipselect                              (mm_interconnect_1_eep_i2c_sda_s1_chipselect),               //                                                 .chipselect
		.i2c_scl_s1_address                                     (mm_interconnect_1_i2c_scl_s1_address),                      //                                       i2c_scl_s1.address
		.i2c_scl_s1_write                                       (mm_interconnect_1_i2c_scl_s1_write),                        //                                                 .write
		.i2c_scl_s1_readdata                                    (mm_interconnect_1_i2c_scl_s1_readdata),                     //                                                 .readdata
		.i2c_scl_s1_writedata                                   (mm_interconnect_1_i2c_scl_s1_writedata),                    //                                                 .writedata
		.i2c_scl_s1_chipselect                                  (mm_interconnect_1_i2c_scl_s1_chipselect),                   //                                                 .chipselect
		.i2c_sda_s1_address                                     (mm_interconnect_1_i2c_sda_s1_address),                      //                                       i2c_sda_s1.address
		.i2c_sda_s1_write                                       (mm_interconnect_1_i2c_sda_s1_write),                        //                                                 .write
		.i2c_sda_s1_readdata                                    (mm_interconnect_1_i2c_sda_s1_readdata),                     //                                                 .readdata
		.i2c_sda_s1_writedata                                   (mm_interconnect_1_i2c_sda_s1_writedata),                    //                                                 .writedata
		.i2c_sda_s1_chipselect                                  (mm_interconnect_1_i2c_sda_s1_chipselect),                   //                                                 .chipselect
		.ir_s1_address                                          (mm_interconnect_1_ir_s1_address),                           //                                            ir_s1.address
		.ir_s1_readdata                                         (mm_interconnect_1_ir_s1_readdata),                          //                                                 .readdata
		.jtag_uart_avalon_jtag_slave_address                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                      jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                 .write
		.jtag_uart_avalon_jtag_slave_read                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                 .read
		.jtag_uart_avalon_jtag_slave_readdata                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                 .readdata
		.jtag_uart_avalon_jtag_slave_writedata                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                 .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                 .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                 .chipselect
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),                          //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                            //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),                         //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),                        //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),                       //                                                 .chipselect
		.lcd_control_slave_address                              (mm_interconnect_1_lcd_control_slave_address),               //                                lcd_control_slave.address
		.lcd_control_slave_write                                (mm_interconnect_1_lcd_control_slave_write),                 //                                                 .write
		.lcd_control_slave_read                                 (mm_interconnect_1_lcd_control_slave_read),                  //                                                 .read
		.lcd_control_slave_readdata                             (mm_interconnect_1_lcd_control_slave_readdata),              //                                                 .readdata
		.lcd_control_slave_writedata                            (mm_interconnect_1_lcd_control_slave_writedata),             //                                                 .writedata
		.lcd_control_slave_begintransfer                        (mm_interconnect_1_lcd_control_slave_begintransfer),         //                                                 .begintransfer
		.ledg_s1_address                                        (mm_interconnect_1_ledg_s1_address),                         //                                          ledg_s1.address
		.ledg_s1_write                                          (mm_interconnect_1_ledg_s1_write),                           //                                                 .write
		.ledg_s1_readdata                                       (mm_interconnect_1_ledg_s1_readdata),                        //                                                 .readdata
		.ledg_s1_writedata                                      (mm_interconnect_1_ledg_s1_writedata),                       //                                                 .writedata
		.ledg_s1_chipselect                                     (mm_interconnect_1_ledg_s1_chipselect),                      //                                                 .chipselect
		.ledr_s1_address                                        (mm_interconnect_1_ledr_s1_address),                         //                                          ledr_s1.address
		.ledr_s1_write                                          (mm_interconnect_1_ledr_s1_write),                           //                                                 .write
		.ledr_s1_readdata                                       (mm_interconnect_1_ledr_s1_readdata),                        //                                                 .readdata
		.ledr_s1_writedata                                      (mm_interconnect_1_ledr_s1_writedata),                       //                                                 .writedata
		.ledr_s1_chipselect                                     (mm_interconnect_1_ledr_s1_chipselect),                      //                                                 .chipselect
		.pll_pll_slave_address                                  (mm_interconnect_1_pll_pll_slave_address),                   //                                    pll_pll_slave.address
		.pll_pll_slave_write                                    (mm_interconnect_1_pll_pll_slave_write),                     //                                                 .write
		.pll_pll_slave_read                                     (mm_interconnect_1_pll_pll_slave_read),                      //                                                 .read
		.pll_pll_slave_readdata                                 (mm_interconnect_1_pll_pll_slave_readdata),                  //                                                 .readdata
		.pll_pll_slave_writedata                                (mm_interconnect_1_pll_pll_slave_writedata),                 //                                                 .writedata
		.rs232_s1_address                                       (mm_interconnect_1_rs232_s1_address),                        //                                         rs232_s1.address
		.rs232_s1_write                                         (mm_interconnect_1_rs232_s1_write),                          //                                                 .write
		.rs232_s1_read                                          (mm_interconnect_1_rs232_s1_read),                           //                                                 .read
		.rs232_s1_readdata                                      (mm_interconnect_1_rs232_s1_readdata),                       //                                                 .readdata
		.rs232_s1_writedata                                     (mm_interconnect_1_rs232_s1_writedata),                      //                                                 .writedata
		.rs232_s1_begintransfer                                 (mm_interconnect_1_rs232_s1_begintransfer),                  //                                                 .begintransfer
		.rs232_s1_chipselect                                    (mm_interconnect_1_rs232_s1_chipselect),                     //                                                 .chipselect
		.sd_clk_s1_address                                      (mm_interconnect_1_sd_clk_s1_address),                       //                                        sd_clk_s1.address
		.sd_clk_s1_write                                        (mm_interconnect_1_sd_clk_s1_write),                         //                                                 .write
		.sd_clk_s1_readdata                                     (mm_interconnect_1_sd_clk_s1_readdata),                      //                                                 .readdata
		.sd_clk_s1_writedata                                    (mm_interconnect_1_sd_clk_s1_writedata),                     //                                                 .writedata
		.sd_clk_s1_chipselect                                   (mm_interconnect_1_sd_clk_s1_chipselect),                    //                                                 .chipselect
		.sd_cmd_s1_address                                      (mm_interconnect_1_sd_cmd_s1_address),                       //                                        sd_cmd_s1.address
		.sd_cmd_s1_write                                        (mm_interconnect_1_sd_cmd_s1_write),                         //                                                 .write
		.sd_cmd_s1_readdata                                     (mm_interconnect_1_sd_cmd_s1_readdata),                      //                                                 .readdata
		.sd_cmd_s1_writedata                                    (mm_interconnect_1_sd_cmd_s1_writedata),                     //                                                 .writedata
		.sd_cmd_s1_chipselect                                   (mm_interconnect_1_sd_cmd_s1_chipselect),                    //                                                 .chipselect
		.sd_dat_s1_address                                      (mm_interconnect_1_sd_dat_s1_address),                       //                                        sd_dat_s1.address
		.sd_dat_s1_write                                        (mm_interconnect_1_sd_dat_s1_write),                         //                                                 .write
		.sd_dat_s1_readdata                                     (mm_interconnect_1_sd_dat_s1_readdata),                      //                                                 .readdata
		.sd_dat_s1_writedata                                    (mm_interconnect_1_sd_dat_s1_writedata),                     //                                                 .writedata
		.sd_dat_s1_chipselect                                   (mm_interconnect_1_sd_dat_s1_chipselect),                    //                                                 .chipselect
		.sd_wp_n_s1_address                                     (mm_interconnect_1_sd_wp_n_s1_address),                      //                                       sd_wp_n_s1.address
		.sd_wp_n_s1_readdata                                    (mm_interconnect_1_sd_wp_n_s1_readdata),                     //                                                 .readdata
		.seg7_avalon_slave_address                              (mm_interconnect_1_seg7_avalon_slave_address),               //                                seg7_avalon_slave.address
		.seg7_avalon_slave_write                                (mm_interconnect_1_seg7_avalon_slave_write),                 //                                                 .write
		.seg7_avalon_slave_read                                 (mm_interconnect_1_seg7_avalon_slave_read),                  //                                                 .read
		.seg7_avalon_slave_readdata                             (mm_interconnect_1_seg7_avalon_slave_readdata),              //                                                 .readdata
		.seg7_avalon_slave_writedata                            (mm_interconnect_1_seg7_avalon_slave_writedata),             //                                                 .writedata
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                           //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                             //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),                          //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),                         //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),                        //                                                 .chipselect
		.sys_clk_timer_s1_address                               (mm_interconnect_1_sys_clk_timer_s1_address),                //                                 sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                                 (mm_interconnect_1_sys_clk_timer_s1_write),                  //                                                 .write
		.sys_clk_timer_s1_readdata                              (mm_interconnect_1_sys_clk_timer_s1_readdata),               //                                                 .readdata
		.sys_clk_timer_s1_writedata                             (mm_interconnect_1_sys_clk_timer_s1_writedata),              //                                                 .writedata
		.sys_clk_timer_s1_chipselect                            (mm_interconnect_1_sys_clk_timer_s1_chipselect),             //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),             //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata),            //                                                 .readdata
		.sysver_0_avalon_slave_0_address                        (mm_interconnect_1_sysver_0_avalon_slave_0_address),         //                          sysver_0_avalon_slave_0.address
		.sysver_0_avalon_slave_0_write                          (mm_interconnect_1_sysver_0_avalon_slave_0_write),           //                                                 .write
		.sysver_0_avalon_slave_0_read                           (mm_interconnect_1_sysver_0_avalon_slave_0_read),            //                                                 .read
		.sysver_0_avalon_slave_0_readdata                       (mm_interconnect_1_sysver_0_avalon_slave_0_readdata),        //                                                 .readdata
		.sysver_0_avalon_slave_0_writedata                      (mm_interconnect_1_sysver_0_avalon_slave_0_writedata),       //                                                 .writedata
		.sysver_0_avalon_slave_0_byteenable                     (mm_interconnect_1_sysver_0_avalon_slave_0_byteenable),      //                                                 .byteenable
		.sysver_0_avalon_slave_0_waitrequest                    (mm_interconnect_1_sysver_0_avalon_slave_0_waitrequest),     //                                                 .waitrequest
		.sysver_0_avalon_slave_0_chipselect                     (mm_interconnect_1_sysver_0_avalon_slave_0_chipselect),      //                                                 .chipselect
		.timer_0_s1_address                                     (mm_interconnect_1_timer_0_s1_address),                      //                                       timer_0_s1.address
		.timer_0_s1_write                                       (mm_interconnect_1_timer_0_s1_write),                        //                                                 .write
		.timer_0_s1_readdata                                    (mm_interconnect_1_timer_0_s1_readdata),                     //                                                 .readdata
		.timer_0_s1_writedata                                   (mm_interconnect_1_timer_0_s1_writedata),                    //                                                 .writedata
		.timer_0_s1_chipselect                                  (mm_interconnect_1_timer_0_s1_chipselect),                   //                                                 .chipselect
		.timer_1_s1_address                                     (mm_interconnect_1_timer_1_s1_address),                      //                                       timer_1_s1.address
		.timer_1_s1_write                                       (mm_interconnect_1_timer_1_s1_write),                        //                                                 .write
		.timer_1_s1_readdata                                    (mm_interconnect_1_timer_1_s1_readdata),                     //                                                 .readdata
		.timer_1_s1_writedata                                   (mm_interconnect_1_timer_1_s1_writedata),                    //                                                 .writedata
		.timer_1_s1_chipselect                                  (mm_interconnect_1_timer_1_s1_chipselect),                   //                                                 .chipselect
		.timer_10_s1_address                                    (mm_interconnect_1_timer_10_s1_address),                     //                                      timer_10_s1.address
		.timer_10_s1_write                                      (mm_interconnect_1_timer_10_s1_write),                       //                                                 .write
		.timer_10_s1_readdata                                   (mm_interconnect_1_timer_10_s1_readdata),                    //                                                 .readdata
		.timer_10_s1_writedata                                  (mm_interconnect_1_timer_10_s1_writedata),                   //                                                 .writedata
		.timer_10_s1_chipselect                                 (mm_interconnect_1_timer_10_s1_chipselect),                  //                                                 .chipselect
		.timer_11_s1_address                                    (mm_interconnect_1_timer_11_s1_address),                     //                                      timer_11_s1.address
		.timer_11_s1_write                                      (mm_interconnect_1_timer_11_s1_write),                       //                                                 .write
		.timer_11_s1_readdata                                   (mm_interconnect_1_timer_11_s1_readdata),                    //                                                 .readdata
		.timer_11_s1_writedata                                  (mm_interconnect_1_timer_11_s1_writedata),                   //                                                 .writedata
		.timer_11_s1_chipselect                                 (mm_interconnect_1_timer_11_s1_chipselect),                  //                                                 .chipselect
		.timer_12_s1_address                                    (mm_interconnect_1_timer_12_s1_address),                     //                                      timer_12_s1.address
		.timer_12_s1_write                                      (mm_interconnect_1_timer_12_s1_write),                       //                                                 .write
		.timer_12_s1_readdata                                   (mm_interconnect_1_timer_12_s1_readdata),                    //                                                 .readdata
		.timer_12_s1_writedata                                  (mm_interconnect_1_timer_12_s1_writedata),                   //                                                 .writedata
		.timer_12_s1_chipselect                                 (mm_interconnect_1_timer_12_s1_chipselect),                  //                                                 .chipselect
		.timer_13_s1_address                                    (mm_interconnect_1_timer_13_s1_address),                     //                                      timer_13_s1.address
		.timer_13_s1_write                                      (mm_interconnect_1_timer_13_s1_write),                       //                                                 .write
		.timer_13_s1_readdata                                   (mm_interconnect_1_timer_13_s1_readdata),                    //                                                 .readdata
		.timer_13_s1_writedata                                  (mm_interconnect_1_timer_13_s1_writedata),                   //                                                 .writedata
		.timer_13_s1_chipselect                                 (mm_interconnect_1_timer_13_s1_chipselect),                  //                                                 .chipselect
		.timer_14_s1_address                                    (mm_interconnect_1_timer_14_s1_address),                     //                                      timer_14_s1.address
		.timer_14_s1_write                                      (mm_interconnect_1_timer_14_s1_write),                       //                                                 .write
		.timer_14_s1_readdata                                   (mm_interconnect_1_timer_14_s1_readdata),                    //                                                 .readdata
		.timer_14_s1_writedata                                  (mm_interconnect_1_timer_14_s1_writedata),                   //                                                 .writedata
		.timer_14_s1_chipselect                                 (mm_interconnect_1_timer_14_s1_chipselect),                  //                                                 .chipselect
		.timer_15_s1_address                                    (mm_interconnect_1_timer_15_s1_address),                     //                                      timer_15_s1.address
		.timer_15_s1_write                                      (mm_interconnect_1_timer_15_s1_write),                       //                                                 .write
		.timer_15_s1_readdata                                   (mm_interconnect_1_timer_15_s1_readdata),                    //                                                 .readdata
		.timer_15_s1_writedata                                  (mm_interconnect_1_timer_15_s1_writedata),                   //                                                 .writedata
		.timer_15_s1_chipselect                                 (mm_interconnect_1_timer_15_s1_chipselect),                  //                                                 .chipselect
		.timer_2_s1_address                                     (mm_interconnect_1_timer_2_s1_address),                      //                                       timer_2_s1.address
		.timer_2_s1_write                                       (mm_interconnect_1_timer_2_s1_write),                        //                                                 .write
		.timer_2_s1_readdata                                    (mm_interconnect_1_timer_2_s1_readdata),                     //                                                 .readdata
		.timer_2_s1_writedata                                   (mm_interconnect_1_timer_2_s1_writedata),                    //                                                 .writedata
		.timer_2_s1_chipselect                                  (mm_interconnect_1_timer_2_s1_chipselect),                   //                                                 .chipselect
		.timer_3_s1_address                                     (mm_interconnect_1_timer_3_s1_address),                      //                                       timer_3_s1.address
		.timer_3_s1_write                                       (mm_interconnect_1_timer_3_s1_write),                        //                                                 .write
		.timer_3_s1_readdata                                    (mm_interconnect_1_timer_3_s1_readdata),                     //                                                 .readdata
		.timer_3_s1_writedata                                   (mm_interconnect_1_timer_3_s1_writedata),                    //                                                 .writedata
		.timer_3_s1_chipselect                                  (mm_interconnect_1_timer_3_s1_chipselect),                   //                                                 .chipselect
		.timer_4_s1_address                                     (mm_interconnect_1_timer_4_s1_address),                      //                                       timer_4_s1.address
		.timer_4_s1_write                                       (mm_interconnect_1_timer_4_s1_write),                        //                                                 .write
		.timer_4_s1_readdata                                    (mm_interconnect_1_timer_4_s1_readdata),                     //                                                 .readdata
		.timer_4_s1_writedata                                   (mm_interconnect_1_timer_4_s1_writedata),                    //                                                 .writedata
		.timer_4_s1_chipselect                                  (mm_interconnect_1_timer_4_s1_chipselect),                   //                                                 .chipselect
		.timer_5_s1_address                                     (mm_interconnect_1_timer_5_s1_address),                      //                                       timer_5_s1.address
		.timer_5_s1_write                                       (mm_interconnect_1_timer_5_s1_write),                        //                                                 .write
		.timer_5_s1_readdata                                    (mm_interconnect_1_timer_5_s1_readdata),                     //                                                 .readdata
		.timer_5_s1_writedata                                   (mm_interconnect_1_timer_5_s1_writedata),                    //                                                 .writedata
		.timer_5_s1_chipselect                                  (mm_interconnect_1_timer_5_s1_chipselect),                   //                                                 .chipselect
		.timer_6_s1_address                                     (mm_interconnect_1_timer_6_s1_address),                      //                                       timer_6_s1.address
		.timer_6_s1_write                                       (mm_interconnect_1_timer_6_s1_write),                        //                                                 .write
		.timer_6_s1_readdata                                    (mm_interconnect_1_timer_6_s1_readdata),                     //                                                 .readdata
		.timer_6_s1_writedata                                   (mm_interconnect_1_timer_6_s1_writedata),                    //                                                 .writedata
		.timer_6_s1_chipselect                                  (mm_interconnect_1_timer_6_s1_chipselect),                   //                                                 .chipselect
		.timer_7_s1_address                                     (mm_interconnect_1_timer_7_s1_address),                      //                                       timer_7_s1.address
		.timer_7_s1_write                                       (mm_interconnect_1_timer_7_s1_write),                        //                                                 .write
		.timer_7_s1_readdata                                    (mm_interconnect_1_timer_7_s1_readdata),                     //                                                 .readdata
		.timer_7_s1_writedata                                   (mm_interconnect_1_timer_7_s1_writedata),                    //                                                 .writedata
		.timer_7_s1_chipselect                                  (mm_interconnect_1_timer_7_s1_chipselect),                   //                                                 .chipselect
		.timer_8_s1_address                                     (mm_interconnect_1_timer_8_s1_address),                      //                                       timer_8_s1.address
		.timer_8_s1_write                                       (mm_interconnect_1_timer_8_s1_write),                        //                                                 .write
		.timer_8_s1_readdata                                    (mm_interconnect_1_timer_8_s1_readdata),                     //                                                 .readdata
		.timer_8_s1_writedata                                   (mm_interconnect_1_timer_8_s1_writedata),                    //                                                 .writedata
		.timer_8_s1_chipselect                                  (mm_interconnect_1_timer_8_s1_chipselect),                   //                                                 .chipselect
		.timer_9_s1_address                                     (mm_interconnect_1_timer_9_s1_address),                      //                                       timer_9_s1.address
		.timer_9_s1_write                                       (mm_interconnect_1_timer_9_s1_write),                        //                                                 .write
		.timer_9_s1_readdata                                    (mm_interconnect_1_timer_9_s1_readdata),                     //                                                 .readdata
		.timer_9_s1_writedata                                   (mm_interconnect_1_timer_9_s1_writedata),                    //                                                 .writedata
		.timer_9_s1_chipselect                                  (mm_interconnect_1_timer_9_s1_chipselect)                    //                                                 .chipselect
	);

	DE2_115_SOPC_irq_mapper irq_mapper (
		.clk            (altpll_sys_clk),                     //        clk.clk
		.reset          (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),           //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),           //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),           //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),           //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),           //  receiver4.irq
		.receiver5_irq  (~irq_mapper_receiver5_irq),          //  receiver5.irq
		.receiver6_irq  (~irq_mapper_receiver6_irq),          //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),           //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),           //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),           //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),          // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),          // receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq),          // receiver12.irq
		.receiver13_irq (irq_mapper_receiver13_irq),          // receiver13.irq
		.receiver14_irq (irq_mapper_receiver14_irq),          // receiver14.irq
		.receiver15_irq (irq_mapper_receiver15_irq),          // receiver15.irq
		.receiver16_irq (irq_mapper_receiver16_irq),          // receiver16.irq
		.receiver17_irq (irq_mapper_receiver17_irq),          // receiver17.irq
		.receiver18_irq (irq_mapper_receiver18_irq),          // receiver18.irq
		.receiver19_irq (irq_mapper_receiver19_irq),          // receiver19.irq
		.receiver20_irq (irq_mapper_receiver20_irq),          // receiver20.irq
		.receiver21_irq (irq_mapper_receiver21_irq),          // receiver21.irq
		.receiver22_irq (irq_mapper_receiver22_irq),          // receiver22.irq
		.receiver23_irq (irq_mapper_receiver23_irq),          // receiver23.irq
		.receiver24_irq (irq_mapper_receiver24_irq),          // receiver24.irq
		.receiver25_irq (irq_mapper_receiver25_irq),          // receiver25.irq
		.receiver26_irq (irq_mapper_receiver26_irq),          // receiver26.irq
		.receiver27_irq (irq_mapper_receiver27_irq),          // receiver27.irq
		.sender_irq     (vic_0_irq_input_irq)                 //     sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver8_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_007 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_007_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver9_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_008 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_008_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver10_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_009 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_009_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver11_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_010 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_010_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver12_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_011 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_011_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver13_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_012 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_012_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver14_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_013 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_013_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver15_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_014 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_014_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver16_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_015 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_015_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver17_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_016 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_016_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver18_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_017 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_017_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver19_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_018 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_018_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver20_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_019 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_019_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver21_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_020 (
		.receiver_clk   (altpll_io_clk),                      //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_020_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver22_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_021 (
		.receiver_clk   (clk_50_clk),                         //       receiver_clk.clk
		.sender_clk     (altpll_sys_clk),                     //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (~irq_synchronizer_021_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver23_irq)           //             sender.irq
	);

	DE2_115_SOPC_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (altpll_sys_clk),                        // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_ready          (tse_receive_ready),                     //     in_0.ready
		.in_0_valid          (tse_receive_valid),                     //         .valid
		.in_0_data           (tse_receive_data),                      //         .data
		.in_0_startofpacket  (tse_receive_startofpacket),             //         .startofpacket
		.in_0_endofpacket    (tse_receive_endofpacket),               //         .endofpacket
		.in_0_empty          (tse_receive_empty),                     //         .empty
		.in_0_error          (tse_receive_error),                     //         .error
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //    out_0.ready
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_data          (avalon_st_adapter_out_0_data),          //         .data
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_io_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (altpll_sys_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
