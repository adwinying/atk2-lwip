��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?�T�RH��'3�g��	4�r�hN�9e�sP;o�k�'�H��2������v�K�]ڥ����R��VJe�_��y;�������m>�w�]g#��e&��>���'Q�*��֬`�9z,��$c���*i��X��x�0�kH!�	��wS�L8��#�O��kGIW��t�.��݃��^R�D���3<�j� �n�M��{8��f`�v��3�?@ʞB+��/�/�1A���_�5(�6��0�,f�2�M.���i�*�&�p�V��8�]U�qb��&6@*�����%�&�Ӭ~F�&y�j��Fv���xg��(<t��WR��-)fM���ϡ�U�j!5"��o�S@h>��xy��y/�����{|�&ճ�/�7��^�˶GY@Y6��6�﹏(�;��{��{�|&qY�O�g�A�rOnk��c>_��%�����X��F���)\i"C�ގ>z_0�^F�������S����4n�hÀ��#g$�#|3Wѥ�FbL~�����rA?b֚��	��]S���t�Ku�n� &Wݰu�b����.�N��̹��I��[�n� �D��v�IM8rZ�e87���:�ІqD�o��_!�KC= ��V�,.@�`:Tҝ+B ӿ?w��C �N�5��#��̣�֢ �q��$0`SɎ�$c�#�i�/���q��>�� g���J&���o;�P�[f��Il('�6+�Ǘ�l��s2$m��OWjdI�܊�G�'up+��(=~Z]�������9?([)�����l��,��<L�g"��Ca�$���=�:Yͻ뼾�0���޼��[�&��c�gH�
�gr�}���C�i��8���o�C��d�O>��w{+��W�(�\Ps;�1�k��p�qޫ �y D�yXf\;?Ё���#�I�����^�'׬��/�w�	d>'�vC�׏c��=�-�����}���B����A3��R7��$[��2U�Y���8�nǘ4��z�6�l���n������pBV�H��.��&+ċ�`&��MwӁ'sW��5�W��^�EP ��G��J�n௣X��ߵ���*�s+���h��G�oIѬL��s�8oUs8,��`��p����JR��~�٤vA<�xH�s��5ܹ���; YZM������=e(���b���>�nʽ��i���6s�&�t!R:���Q��a���8[�t�D�����9�c�׶(Ƣ�+�l����\�rp�cV|�'_�n%v�\�V: ��ބV������2���1���>uܴ�F�s`���h�nG5�xĭ��<��\3p�/-F\'Q�i4�(z}㻳�8�;���X�D.` ��'g��TX��Q���g��8�,dݎ��Hg�[��mٓ�m���N��fdF�Eۈ���i3:���{�
������s���
�3l����mv���I�=Tgx�spj�O����R�dמWi~�U��x2�2 ���@�K�2�?W�����"}!!��k�Yk}T&<��f����w��b�e���<��)���������5Y]�l���咾n^��Z9ѥǂ��R(��F{�Y'-�.��̡����N龨�6U��W�r�m��˛,�ay-a�-��S�j�h<qz��z6{�ӾBﹻ�D���n����O�I��`��
^�$u?js�rpd9��P���sr�pr�FϮ��ID��FlU���p?_�ڈ,�O�s��y ��Ɖ�/�f��	i��G�Rp7��S��Br{Z�,^��?!ߝ�¿*����sClD�QL�X�/YRR��x^Ɨ�z��4��V@�Y���s�d��N�8."b�*k�CH��� h5��_�SN$D��O:Nj:]\�� qsS���+%��\���_,�y�����l�$���/xEܣ�-�2Q������W�|�.�2�vn�43���!��"�A�vg����ʖeKa�@>�S�E߸��n��a�`��?.�_S��۽&P�B���Aa ]���`�o�M��M����R�K̏��2��*�����|���WG:�^qD�/� r���3A\���Vbk���$*���`%W�K�Π�.��B.W@��&X�w�ULc�0�U`��B�X�JjnE���$�v�37�E�H����e���\6����8{ܪt��.�8�Ui�(��}����;���Oz�/�O��u�ۢF\Y���X�&���I&��ek/bZ�+��R&��Ɂ&	B��тx�E{*�5GJ�J���	��&I�������O� :�n4��S�|�3ҼkC�?GW�3�5����/�^�S�$(��F嬃��<Ӄw8r2R�_��`��8_�URh��Q���t��7J��2Ws.���v�|�x�7IP_b���X�5�- Ym�{�C��/z-e!.5����32�Ar��o�p�/����)9G�m ,��zT����7'=���
��5>�ֲf��	��x#�vm�偷z<�k�cq�������a�R�<5R`��SP-�DzC�{�x�:��z�  �Bq����iz��+;���UΈԓ1�y�u��}Y��xzl�|�1�qb��#e����Mt�����c�QU�r
<Q�Յu�F�^3x�B�͓wy��He���q�݅�_ʭA(g�Ɵ�4�b�0�)�Z=@G���i��@��b&G ҄J�zC��9�����=m Qk��_��JR��a��"���Q>�?*����.ګ�i��޶��{�:󽟻�[W"���S,>��,l���&(�
�"�j� 	��x��r�D)��� ���5�l��
y�P�;}*,і�2��j4�=�����<��l`m����([XF���u&���K�?�q�o,g�
��*B�4�J|�k5�oX෉9��F�,��q�5Ҹ�/K]�N#�ny��Ke������E)�P�yrBH�QW�C-��À0Ś*�kã+\JB08��:�������Ͱ		ln��M�W��v𗶓��</�����-1��@���9LVQf↮�`���57�Ѣ�b��9Ue`�bJ�oT��/�^�*�ħ�� ����x�!��0���aڶ��ܝ�2�Ѵ�5J�C���0Q-%���΀���[uחā��C�����|�.�N:�m/(���*z
Z���S����a(����ZҼ?����P)�E��OW��q�0\��3u�l �Vw�P�yt&��k �V�7#�.�v������@������65I���f������i��yۚ�2���<���QD��LHj�K��1��Z-:�����p��_�t���|?2:���͜��#1݉KI�l�DI�����'�y�0�,|4v!~�*N��Wln��Hr�l^�_m�jܓť�z��E5�!��!5M����i}�h�nbM�>M�ZS���8����#X~�!h_쪵��J�����^Y��9�֔L�a��(ӏ����mS�']g��4)Ċdk�N���m�����ˏ�Ţ<�ddi�=���n(�ӍC��^�#���`p����^��8���������H�n=� J#�/O��Ő�sy��Nnx��r�j�o��R��'�{r|H
���Ɩ|4� ���_1Ȯ���o*�u$J��ma�U��ǝD~���h&{$�kG�4�w����	4�J1^Ms��E��9��n�/�|���*	��mx�ά��h޵<I��`�B�f�U�Z�A�ܮ��l���6���7�˝Vͦ�aaJ�SΔ��J(�5��S_粪 ��[o�gυ` �B�}(��s6B�WV(Ҫ�ꁮ����r{6���+�i�`0�X{����xnv��ۖz����)�������Ӥ8b̹۔]vQ�r���ʸ6l�a�H��I{x���*��e�(~�	ۈ�?~���1�	qG�1� W|�CἜR��_Ir�"�3��)ل��AJ_�%N��H�W���|���	#h�=0�)���̹'^zw����3�k߿t�X��P����&o���s_ۨ��Q3}�!1��+ ��r8�QB�[ܭ>Z�c����۫pT1[X�}No%3��Q�,f�2�tjJL�"�:}���BK��D�>���[E���
n��{�񤟯�m�}ow�^no]���.>=�fY�� �R?���$tj��.H��*�G�,�:�q��nX�Pl����5�¯	�R�,1�ѥ��յe�d�VIz������j�(m�iF$J�K����d$���sە,�r|~]�J2�]I�&�|�wM�����}J{'d8�~�I�`jI����wqi���p����m+��������KAl;�G�Q��QO �^���u���lt)�:�y��`Ľ��� e�ϱe n�x����
 _p�;wAH�`2�ۛ慆r7��H'8���d�?��}'�-����G� �����#_�������[�1���=�f��8ӑ��Hw�w�7t����V_I*tS�U}���B��Z��x�\��ث�X���A���NӎS�o��&���5E��+�qJ6=������I
6h)x͚�ɸq�Z���Y�(�A>�k�Ly�bQ# {.�|&����E���\;��]I�/wɪ���~!�`���O��&H6����j�Rz���N��@N�O���k?$�i1c�w
dr�	_������9�S��7��au�f3�͗դg�#�Q�T�1��lN�����+S)n�^\����+��1��e:3I�͜���7����Vk*R���]kS���a3k�>:��Z�Z�&5�~�W*�Q��>�Ռ�MT|��U�\�gzh�-q�Y��=��Z��(����,��>���ocܹ�"T �mѝps����!�/k�S	��<�|�<�^�d��v+''��4\CM&bB?��Q|gTgIUm>S��j��O�ԶuŜT�� c+����ź����%O��4���Ax !�X!�Ɗ�����$�Ď�>��y��y:4�吂v�(�3�d/�A����$kV��/�_�o�T��.�%j���X~��TM��f�s�ϋ�0��K�/H'�>X��%i�W<؎Q���81�v����q���S�t�~�\,xu��Gzt���HKi�t0|��'��]���f�"bq���{\�j	�KX�Ж���z��ezm����&����28���[�� ���/�~�<���Þ&�:��T`�t{��p�~�4 �|� S"i�{<�ӝP!!y���s�p�tg:=�i7��F.�!���N �e��ڄ=B:�R7n��� #��tq�HT��ʢ�F?EǪ$i�L�RF(0M���u}A�t0P�;��r��sHԛn�P��Ɣ��g���zJ�c>	 Xc�sr��\�a���7M�Kb��&������A�
Ga� �%~�=�i�f=)0�����9^p�n>��R�
4įʄR0�:dg��ڌ71?�F���
��q���w���k�(:mG&�v0�v�V��h�n�{��׵�������#��%/��*� p�G������a���S���E�Xa���X�%�-"�[�-�A���%��b�^�hp�����-'��U�#U��t��RS�@{�$�4���mϔ���eG
�/�R:a��qZaJ�B�5]j�
Z�M�7���L�M֙�!�h��Y>�^��i_��5��Uシ}��~�T�:{y���a�-ڃ���'L�A�n��_ �8��|��L<�88�pa�b��5=���h1û�}�3��)r����>x������'���I����<!�?�V��i6���tCvW| =�炑��M�K�K�rb������8Q��ҏ��W����	m��r������d���ǈ�>��>ċ�˟�,�To�ao+y��S�	���#�RIL������wBd�#���d�&���w�S�D�%y���T���i1]ug�\=Mj�]]q�F����>66%K�I���.C=�?�MP���& 8�����V�i�T~�Xhi~2��m���u�!G"��57��U?��K1w\�q�Y�a���*��mbi;�������[|6�W���Q�U�8� �����ꨋ"	8n�0p�m�"@�����`����z�ȡ	�`4,�� #�cr���mww0s����